PK   IqwTq�3B�  7f    cirkitFile.json�]]��8��+ϫe�K_�ػ;@?�t0��}Hɖ:�8v���tO�������E�L�&l
�q�&����.y-����X�V���X������_��x��P7���w�r���C��|����l���x���X����i�W��T�����Pq�gyŲ�DYei�n
V������|NF`'s0"[�A����
I�@E`�"sPW�r}��x���s!T]�*QQU�*RU���2�*�b&��<�"���d�15s�!$�C�"�"%s�"�"#s�F"1K37bU1�#Us�I�D�Ȫ��J7Rg$��L����2}p Ch��
�Y�3<B���x2�fA��d͂����=ߒ!4z�%Ch��K��,詓��qz�$Ch��I��, �cz���I��,蹓�Y�s'B���N2�fAϝd���������U���Ur�&��;p�v9Q����H_/�U��8�x�T�c��y��S<v�q{�Cw>!����D8�eǱ��L��jeǱ��5��N`����Xv��X�$V;(;�e�
��Na����Xv�����X��8�+�v	V;(;�eǊ�]��ʎcٱ"�j�a����Xv�ȱ��X��8���w ��+,?�g�z��CW��\_pp�����3w�����,?�g�WX~������6��8���/	�\q`�q0?sG������`~�^0X?p������]l�~��ˏ�����������3+����,?�g�<��C��@�� �\p�������:�~��ˏ���2`�����3k{����,?�gV%���X~�Ϭ���?��8��YS�\`���.քI���Mɸ�DJ&IT����4-�D��Z�֖��݇+n'v.���}��ub���ԉ݇�J'v.��}��sb��RƉ݇����5�qg�o�ڟy֞�����g��ڟ}�މ����g�W�ڟ����g��ڟ֊�����g�b�ڟ�j�1�$1�$u�%Ɵ$Ɵ$Ɵ$Ɵ|#�|V�q��v��6\[L�r�p�5VYʳ�,��Jrݹ�Q�4<qR�&�DU��6��{?��	�}l�]����DԤ"�TR��l����Z����`���}Ѝ��3��;nO�����7{�)��ǎ��T�y|H��>>"xu<�'�D<7�JL�N"��@_)_�o7F=���p��,��ڿ�g��z@�m�Q�4��2(F �֓��:�`�@�f�ih�b�(׌���(A1��:F ��_è�պ�4F9��3��H\�ƥmRg������QH������q!u�< N��a)����8��:�'X�<�B�}@�`y\�&�<.`y�ԙ �8���qRg�����QH�y���=�S���x�ds����Qە#T���
�j��Q����j��`�ц�u��v��(0\�G����Q`���
�5W�q��p�7�k��F��p8*P�\m��õ�pT��!��.>�k��@]Cp�~0
ג�Q����j���f�a
.�k4�Sra�0��"�Tv���,s<,R�0�W�c!<,R�0�W��!<,R�0%X�C"<,R�0eX��"<,R�0�X�##<,R�0�X��#<,R�0%Y�$<,R�0eY�s$<,��B��,[�q�m��,[���m�[ba�2����6L]��Ì	��6L]��è	��6L]����	��6L]����	��6L]����	��6L]���
��6L]��v�i ed-�t) ��z��R ��5��� (#�~��MPF��ΰ�B�`�wl�?*&��vG�0�B�`bxl���*D��D��~�vVL�m4��q���D����WLKLKLK�T�����v{�gP���v�O��2���	��P����[T]�F��o��Q%fL�~�|��>G��Lo����۱��@��b|��ގ_��� _/���WS�ӹ<� S�}�t>��K~�L� @����35�0u�FF ����ԙA��:S##Pgja�L� �@@����75¤H\�ƥmX��čB�M�0�`��Ò7
�75�p��oK�(����	��9,���zS#'X�<�B�M�0�p�o���,���zS#'X�<�B�M�0�`y\��8
�75�p��q��cH S#4j����05B�¸:L�Ш@]Cpu�A�VE�Q�����05�(`��F�u��ajQ�Z�F���������
�5W��Dk4�k�S#��
h4*P�\�F���hT��!�:L� 
X+�Ѩ@]Cpu�af�a
.�&3�Sra�25��"�Tv���l� 8,R�0�W�.S#8,R�0�W�.S#8,R�0%X�.S#8,R�0eX�.S#8,R�0�X�.S#8,R�0�X�.S#8,R�0%Y�.S#8,R�0eY�.S#8,��B��,[���m��,[���m�[ba�2�&��6L]������6L]������6L]������6L]������6L]������6L]������6L]��v��ed-�S#:��z��Ft��5�3L��(#�~g��QF���15�`�wl�S# &��vG�15�`bxl��S#@��D��~�9�F L�m4�cj��D���9�F LKLKLK�T�����v���QnG����v����QnF�����9�65��`�܌oS#:��x�65���T������R����b}���v���._.>m���xܕ�zSl��ḩ�����_�s��������aI `�d���'*09�?#��3�]}�����G�ٓ7e��|3�ō~�3څ&0y�A��)5:t��%�U�9D~[��ǽc�������5��4u���_��~�������o}��_���&/�^�^���ur��~z��X5·x�F'��34�n!�&��Q��	��?E���z��[�����a��x��B
��N�!�������kΟ$"��uO���s#^�}h��<T�i�<R���JD��1D�]�Q�tRd���Dd��D�>A	�TL'ۤ�EUB'E��AdA��Ad��'��H�tRd���Ԕ�ȼ��K���@�H��o��c�<����<����< ��2+�l��T� �
@>�c�d�� �S���� �S:F��*@>�|J���@�ȧ�O�����c�*�\��R��x���JI�s<8���xX�������\Upx����@ �圂Ã���x��x-wD?,?�#��k9��� �a�9]@<^���������ZN&8<�~X~�G��r+��A���s<r�x��#	�������.� ���3^t	f�zx �!�A�!��>�!�3t= ��]���L����%	������]���L���ѥ	��ˬ��]���L����%
���|��]���L����_��u
���L��]���L��L�u�m7�h��S�]&�@@���:��ev�h��S�]��@@���:��e^�h��S�]&�@@���:��eF�h��Sn0�a:O�o�V�a4O�o��a.O�o�Ɯa(O�o�~�a"O�o�'�cO�F��qd�M<	����9��$ j���X��25��s�I �H��ϱw'P#�^>�̝@�DI�DI�DI���(��(��(��(ߊD_CvJǮx�!���Fv�����s1å} '	p�����m���Dx������ߙ��t�;Xoo�����՝���L����Jޖ�~׍��� .1&�0ۍq��'c7��w��M�1�db�D��ilR�?�Yc,cx�д�)7m�i�Mkn�sӞ�����h�Maz�C����Gk����H�C���czH�C������A��H��|��W ��'���`���	������SwB��ٜ�B7�PV��}SN�H@����=fR����۩���y��Î��W���G������ٖ�27��O�	�"zj�&��ytɮ���}v�[��>���;�q�#�$�d���?R�G��(�?�폒��v�.w��B��9���l���,�(��4^K�k�DK�Hjid�7Z�M��tP����/����ٌզ�n��Pn�)B_:�4��<��ʅY�%����S]�y��Z�B1V<=�q���J��"�W��_Z�I�؁��%�N�U�K��}����X���L�쏇���=�u��'+��y%K��U��,I{52l��Ǎ>u%�,�F_q���FGn��בX'US5q�f��Mϴ��~���,��V3/;b�����d�������}���x����ɇ�{%�*��g,�D���v<O{����J1�	ս�6�J�"{�t.eN�T^�k�8�*~0S�<KT�=_(#pY��%IOD�<}��ܞ>?m��_��S�����+����L&�8e�4��˔�x�I�˄_��uRעn�h�**+�#}F���&�!�E�&���5A���b�>�Y��E�2'BK�x?Q���/�B�Rj��qo^��떧�q��U�ڗͿͧ��o�����?�q�'&�=��J]��:}8|�i��yqט�?<��_��m��_�;��z�k��Y_��},�OM�>?��4�)\6{���cy��_�� *�ђ�l�/�����1��sh_�2׺Jj�z]%e�&�:"�,�X�5,�׼��Or��yř������-��\6rs"��T_?J�����F5R��D���WL��x�I�͆�eUn̥oeA��s�H?�]"�X��!`)3���$v}��RƑ�fRy5�~h�M�Σ�����}�"��ک^:�Nݑv��[��H����.��¦��k��4S�pB���ã�� �|o�
��H��ڐv��hG+G@;Z9�����v�.�ﻂ���ˎf�Pi6��f�@v7��x��0��f���)���LZq;�l��Vèu��,`��3ꕐO�22�2=�N�g�W�撪������ڇ�*�Re�]�dU"�YU����<�eilN̰"23�4IG>ɒxϻz� M7�-�Mux�o������>�HOnWJO
������~8_��m��`�*���G���n�w��*���~��kl�r��Po~x�������_����5Q3����E�X������/y�˧�~���S��x~����i?"�0����n��-Ա���Mz�驊�����g���q}<l��w��C�����~a
韚w惟�	�ɼ{���z9�+buq���?��魺��j�tA��q�D<��)�VWE���×�������껃nv<cV�ގ;RL�9Q(D�:B�ؠ�H�&7}����W~77��+ᛯ&p�)^�h�(�����J]�z���j]rp��p��^�[�eUZBrxں+���z�=:bMi����`\�Z���i�tX�tSo�"N܊�Y�PA&f͝���:�6/?��W�^s�ݭF���{�p�[�^'��ί�	�@��O`7�_��(�od���l0M�k�����}[]�Hߘ��>�D����3�Y�P�3k�&��|��6�n� D�xV��9��$"�̄,|f�İ��ʚ�h�g3���j��"��\C�2`ᓁ���j�'W��^n۫�V�I����)~���F
�D�5K�o\��8�)�V��/�k�8�75�[/n�Q���	T��J�<��jY�g+�܁"�&�k5N��v����[y���rg�T�;���������?��<�O��,��PK   IqwT�Ʈ�"^ /_ /   images/5007451c-e503-410b-b74d-3a3f8b63c8be.pngtwu\�_�/�HJH7��4�0�
� �"Cݥ� !�R*)C7C()]�1�0��y�s���{�~��k�ܱ���+VW[�>)3)�}�W/^������	#����S$��ow�뵪2^�(��߁.�D�^K��/M����?*?�G���A����������4�?��y�I�	�G"��/�h`�m��)kq����	�����+yٿ�+�ۆ�����K�_��h����a�<��og��&Z���!� NIaQaч������v���_�����Hᡃ����������@�	�����!���m�/����_N����������#č��[����Ç���W�W ���Er�����.P��������f��h��1�G�/3�����Ǚ���?���+������ y��U�?-�C\ ���6� E���7���俼IIK��8&�k��-�������l�?���n������ȿ�P�T^���"���/<�gxj/����yY�|�Jȫ��� 4�r�}�"�������[4�}6��,t�����J}�B_=�
�P7LQ�i�b�|�0O��]�e��k��1sHHH�������r�X��֒V�j���9��A_yºWv[Z��Y��o�p��[4�͈Պ>��di�"�Mo��\�u�h=6�լij���CU���F}Z�"-d�P�	5�U^��0����y �i��Drΐ�LcL�;�֮B��7{{����Mp�5���S\��7�`���h�[']��X܎"1n�^�������SMZGB�O�j�}�\;~�8�8�a8?:�Ǣ��UV�4��m���ڨ^�5yB���T�zو��J}D:3��98yR^�n�i.{�1ɝ�V��LHq���AYOL��̭�����u�q��.�O%�N���\�8�v�K����%�)�80����h��D-�l6؅5�lCr��eW[1}[!�I��i"SP�l�r��ϝa��}���?!T��������:������m.T�������{(�S�o	�wڈ}�.6@��Y6ҧ	��`����}�/�#�jX�oTH�~l���b�)p����C�m�_~/#�!a���K���ږ��*�sI�f���w�7!��d�9�FtQ@��7�����z�닂\����q�#���.]�lZ��������I���a2X�b\MM�D��C@��g�~���s>�uc�^|oo���'s�M�ޞ3�KJ�t��_�Z�� L60�Tհ�k&~�v��r�{�X� ��G~�L"G���pu�:��ǀ���r�����J����oU^����I���:=������?��\`@���#�,^��ȷ�HFL� $��DH���@����N���X�s�SbQe��Yʄ�����[���G��.��h���)ڵ��Α�M�Qk�6�:�	�	�����g	`���F��,e�6z��	;�Nh�{�x1���Z��
b>C/�Y��uۺ�wKI��L&����B��/d��[0�+F,X1"�N`mQȏb�+�"���\��D:� r����Őq]}�Y���O7�����8��[v�k�3�Z�����H��TXe�)?y��ao©��|hC:�!m�G�@�*��\�l^(�,n;��f�׷\���X�db΀����L�5���H�%����K�il�N*�cwRC����<��9�Z��9ΐ%��]B����3Wi��H�~`B7�+(�f�ì�^r�+I�5�`��oWN:`��� V�L�z˘�������X�wU���S�^]�q5�h�;pR[U��3m��!	֧:QϾ�X��.]�6��a�| �?�V�t��O�Ii��}Y��NÁG��[H�����Ik���b�������݁�d�F�����TTT�n�L--������iL�y�x���*&%&޻螎5d�%("h/�G9'\���yJN�q�/�D���>�,=����by#)�+��������܎��L�+�ϥ]�gñ-�7�tq.���?���2=*�X���tU�0X�p��	aUl�fZ�B��>�E�4M�WfY¢.r�Ns=�Lq�)5�%aK�@����DG_U8�±�7$�(WV8���V'��Ǚ�-�6�|-����6�A��=E!n��C5ղ8~�6�vJ
�'�`쟦P���秃�Q�����w_?��Z��d�����
k9}ꊄ�y���y���QF�8^�f8ܛ�el��"i���G� �|{�W��+T������h�����0�ř���ג\w�O6���F��%*V��_,��现9��D�نil�T
�s�$Z���,T���Fu}=3f�"�����jc�m�gʢ�3$1=J�O!�N������;�����ҍ��1D�ɷu���ҳ��l��L����Yf�F;��^��vc�1\7hW"�����ߟ�/�*�N�ە�߿{_�1��ZS��<�Y��w����sb�<��m��\����X�u0���#�@{��{s0V>�b�*Y���,Kx=\1����7��-��n?�שE%��]�����OW��$��4�M2��	�L(�gi[_T,Y�ܧ�H�/�k0��˭����v��-�*�$ZG��I��ң���ɯ�cb�GJ��|&�i�4��O�N"I�x^&����u��K��{F|�v��\��^�E��?����U�ϩ7���cH���q���2]�>����/J_	�SN���5�F�P�s��^���Vů��OL:�\���-	�_�`G�ܴ|��
�}��3����?�S��]���l�l8M�`X�hP�|+�����p�c����ŭ�v����������NM����)dw��0�:_2���k��R%�&}�L�����u�����쥀6�N�]��N��b�g̾�`�䍃Q��>I����P���96+v���ײs挋J����Uj�P��d�'��-�I�˽r*���܃�C�F�O��f�����rd��,��W��]���m�f՟k��RR�.�h��[{�i#��k��Q���8g����t�� ?}�U�#��J	��@1.�W��ISC��ι��6W�o;\���cff�s�\:_���>�v�e[�t�Z�zD��6m�\�����?Y��d6�sw�*ww�ٙ�eֱ9�ٕ�{� ����\�Ue��Ϭ���4qiy�F�&K��(��\�ӟ��L�t)����K�G��20���>�����V��b��3��H�-2R���� .��W)fU�a�� &p8�ݘ�&�E���"o�5�aiww��x�
�_R]�{�� (l�� )�y�bit,�P��4��	�B҃�&���w�g. ������]�q�`���b�Dl��f��X�f�k�Թ_�� ����5_T��F��͜�\�w�vX��⽸(�X�阀���넌 F^K��l�!�tW��gG� $���$$�#xԛD�rC�'4�w0I����4��dg�޾:DU�>�|�ڳ����R<�F�m�Z��}�3��mY��5�+P?�7�=����Wf���*���r1�s��`���N�:q�����;5뎧�hqƧ�[��)K�G��܀�����J���̞�i�9@;}l����;.y<P�\n[��B���պ�8��I2�	�1[epE��@��v-����V:F"uJ���p9*9�����f��ֻ���zLNP�*f��`s���x��s�\t�cD���6){��˅|�P�at��v4�Jgܞ�嬠gz���O�mh[D�S}hq	�2�m����~����5���1�؂������?-��}t�#q��>��X��c��,QJîB7M�'siE���j�9+ �EZl�9�<�DA��ϑ��'�g�g���;�<@Sc�����ɯ���dGU�`V�q���<�p�eF�M����N9�����F���Q��⚐����̱����̖�QSS��)3��#f?ɵ���#Z�S�;^$���RI
N�}D��y�V >�js��y�Ⱥ�ܷ�^Jp6�"��^��,�H-�P��j.�����,��`:I����R��(��1j��8`w}ڈ�M�ʃ�&�0�4XR��?UX� )H<�M	5�X�2���r�>�0N,� ��\}���]P��x�/����U�G�uu�Ns桡��kD6��L�h0.�Ҿ��w/����(�wB`��9��X�ٮ4T��mۤ�H�l��K�|�ߥ�eq�ߡ���S�i�t�NN�zͨ�Zp�eM�n�gD <��{�:3c��ngupw�7kS�2�� t,WA��7C�j}�`o�|�c��yl��@C�����w�Z��sQ���q�'�b�� T�)Q47�9ʍ+��}E
<�x'�j�2hfn,����~4\�&�h���ur����;MMW�Y�LG������Dc��U?�O��'d�[�.�Ԥ�4��KZ)�[ˍJ�$ێ�b?n�A�+� ݗ����MK�P?Ԕ��1]��ꖗ���G|jef@r��=i�oar4ň<�u��nM�%K']��tQ`��#����� ���,mm_��Z؈�����9��@��w��S�Y��EN�ɀp�� �{���wP9�k0Gl���+��I�cw)������ߺ��w
@��gH�J�Õ݋��Pk����z���My�RRRz������&��#X'�g�xי%^ӥ�K%���W�6��LÝ:����猌,4� :%�S˨��s��.����H>.j��g�#K�sg�i�`D�u
ow2SÄ��҈�yT<Ĥ������J�Jǻ�G�ke�R��RCz�]c�:ٞJ(�ʴi�T�q����l�`?�N���3QQ�R�!S��������p���?>>!=d%��w�g�ES��VHZ��D�F6�IS{'�t"V'(�!��9]x:
0x峖e3ۿ�g�H�t<p�����/�c�ar��ɣL҅�@�z��!Wi)�I��磌D��t�i]ge����P�� %�����Dvf��o�`�^�US'���B�Vd��1���Tv�aq<=�=>R�"	�n��2.sޓt�;|G�6Ƿ4��g��"Z�N~�F��׸�	{���Ml������7���B"i�I����i��ԃ|z�͌[Ѻq�DD�~*�ֆҜA�w�l<>ٞ�d��	��Җ ��4�<Y zS �r�|*m ��TbvI�P��a_h>=�e�b�+·!�\�2VYo�]#��?�=Zf��=t���!���-/�i�D+	�ފ�0v��B�������P>��q!��&ѐ�A�NK���W��>�F�b�a$:=��,���xEo(L�}˯o���1� �t�[yC�PQ�paa,ӌ 2�#r�k�<���������z� }մ�^���CL���C2�cN�=��Im��I��x��V+&|�J��UR��d�(\��l�ɑ�mVԣe��N��b�חb�����t^������¢�>��g���/��L�K͈~2 m��L<�{_z9m���QU�j=�hЩ¥�� 1��ui��h�P}u��=����hoK�(T���߬J~�:���{����ʖ��G�zdT4�-�6N�D�q��<�ŃȪ��+i�Io��S\�y��B��GK)��$��S�׉�����ǣ��Bq�M�}�aϬ�z�Y�x�mŃw%���aRVT��&:]uI�%B�K!|��(s�TE�� ��=8�󡥷���n�U[����*���i�+��R_,6����s�3֞X
�4����j���P�Ч���
��йl���  `�^N򞩰$�R�����v�<Z�-h=�E��������Yɮ3J�`wi�{�T]��w�
j1�k��M���bnB���3��ͥ�_����0g5�������q;ٕ���r������>�!��r@E��K�����^2�|�%�I�bu jA��\.��`�{��^��	��j��ӎ�)%��5��A{��{[-6'�ks�D�ޠ�p����TG��F�åV��YAD��6$}]51#4r�㲥�t��B�2{�r�r&d�L����e�uv��l 7{�j�l������@���3+]�+w�>�qGN�$۪"�*ۭ����߻�=��7���FH^�(��a�����^*D�?ߧ���~��U�?�gqx��=���)_m��]����o���L�t1xz�o紺_��I��V�6`,�㸿T��<���e�y<�������cԻR���q��מ�����7�r��i�E7[��T�rd,��(�#oU��Ѳ�8U�0���z]�c�f�T�Ë|�����R7����]&�U�n����� ���7��vж�e��x}�+83�#Q�$�l^�$t	����~��a8Q��L	��6\3�ƭ30�����ǚ��
��
݁�,����� ,��V�V;��ݻ\5\R^�:TX��qׄW�C�����,�3�p����A������N�+N�f�����2�C\���L��_�����,��sDl�zV+7uU�#J "6��`9N{�3$RbM(tt���I��a�e�H�F�D_�]V�S�n�l�j��t���}�=��!yq��|�yM��ka�GOA/7��J��kν�E��+ݍ��||P���ݐ��l���M#��|VZ����H�?ߋ�M�v{��[+�� _,b��T&5쿉��g]W�SE&����k�2�~��`�;M�V�M��r�#���
���e1��K�gu�XB�!��SnY��f���C§h�Wt���H{b�Β���X��x\��RP��d�ŃN׏��tX�R|����xT�����s=� �i�|o:�5���ty�+�^,�Ս�HF��ei���'���ܬ8Da�����B����<xg��e�=��FL~��B�z���6������z����!:�S���9_*�G�)��QW�hB�5[6F^���'��Xޅ2 Ҷ��(P��ТG/���~|��l<U�1�cڏLs���Z��L�V��Y�
��j2W^���YI2z��m1��5��o�kD�p�8)�}��V��K��* �$Ayv"��'��b����D�W�<�<}���u�O*.v��7N��j9���S���@���C��
I]^Oi�N	��;�O)�<�2�Rӯ��l�=贋eu�+}HƎ$G/ ��{��]�u��*ʲ�J���D��٘�Y����i2�Eٓ�M%��w��i��ۙe�f(SIx~�ds��F���L��i��`��m��m�+»�ɕUĲ�4W�oyz�c5�?ԭ��C�3�����Mf�}��ZM��{����>Z�o��*���Wޙ1*3�G���,�g��d���=pC�<�ˋ��bҧ����5'�{�}%C�{\����� Y<j��AML���b����q^b�	q�v�%i�-u�f�\(�z"|*Y�r�T��=w�0�Z]�!���G���[^d�9�]� ���={��mF��$�5��Մp:1&�4��GT�X��AT7Z<�ox�����n��FRbtµ�~4��i�t�0Je2u>vr�iZh?���ި�� ƭ���i�vgư��ۅ�>�J4@�sEJ]ȽV,l�N����L*��l�lGRb8ћ�*
���9R@pf�#]��3Z�nOs�T����V?o���P�}��-�p�A�L�o�w��f��*8뺞(��Rtp�H �ǫ����k"��p�|.b���s�%Ck]N�=�I�ͤd�2����6|zkv�4���/��P����ǈV'�CN�rDE9�='$J�+'�LS����g����Ro�Ɏ��om'~�=j�޹��[�R
������n���1�g��|d�m��N""�	�
H}�N�+�%�|G�DJ�������ȍ�	�u7�ƕ�@�B�,;����de��{�$Nt_[1�l)d�y�S�"/~�擔��R4ݥ�����*`��S��z� D	�w�<W�r9�#92���ȼtH�^K�HRw=m!��R?tc{��dO��#����F���f=�+�� u�*� ��+eM����T�韙�.s[�0��[�K������ ���U���W����v�~�Yz��h������ަ���[�����d{�6��5�e:~ܮ�����&����E\�)��Y�xڮ�����iYhb��W�3����N��td�2S��EoN�'nz���G@\O>A�����r]�����*�G�+�@&ˋ���Q5�_1{�ZY[|I�$��}Tf�JL�eW�޶_���g��߷=����D�Y��|_8�Ꝗ;X�90����q��@ OZ�\1���
�P"�'�3���A�Nj�D��;4��D��QӦ�yE!sS�%��PmV�bJM���cT��B�_�"�����+gM��6��y�. ��mG}��(I��s?;J^���U?�D��`ub�k	�ڕ	�"=�S6k.��ԯ4)=�4{��JF��P�cY�̿��>iǍ��b�����d��L1�Ǒt�E�1�����P���"�N-mp��\�c��Z�Ԗ�.��4j.+H)���u"��3"���%�8��|��Yj��*����Z��{ih�:���1x�JF8ZӋ�[s�ّ�]W[!Ε��!��lK�Dg�R��7g?���D���[��my�IS�!7� U3��Z�$�����]�w���{��n��0[CT�`���+�cG�<��-�_�\���q1���E��^���Qa�8�t�H|�]�
�K/Wt,�o2*���1O�^�<a-�E��CE_���=]�0ۋ��'K˔i�y�&�R�U$����P#���&t����yH:�w��"Mɖ��e~_���l�OG�9��?Y:pg��B�2HY.	i�q����^�Q�b�)*�Dwb�,'�� �V4/�F��oE����Fy��a扠�<��PCc�qZ�zmW��-){�����$K���dWUi�ZG)W���!��O�*�D���Hݵ��V1��}�G�s��!���U�'�$6t��so�N�����ah|TQͮ@������e�0�w�2_MD�_�Ql�j�=����xs����T+��'j�u��׍h˹��qip�� |롒W�E�>��oE��e���67�㴋:������.?������ ����#�GY��h�Q �^��\pijR�3���3> ��2��Ư<N�3Ɠ��
�NW�\+����D=��b+��F��8έP�o��Z�J�`Rm�t	����c�Iug�5
���˦��ҫ��[O�̄p�~7�`�u�p|j�:��ײ1�/k[��z�ʴ�g���O�&�j�&��*`�@j������e���w��TCZ�c�ֽ�g���2���bfaI
*�4�IU�:����ƴ|3�J���R�[v�׊�&ǐ�R����%��Fux��w�$��A�%�j������}:���}�h
�~L^??iD\�&-�p� ���4~+�p��yn�@�����aw5��>J�z�	�)Iu����9S���xV/�W3W��"��N9y�U�=|���S��m?�(\DU�n�-��O' ��W�6#�,q�g$f9��%��Ahrx�D�aft�k�Y���8��u�n��p�8aج�bX�����b�?tD�8 ��2e����~�(
B�.���G������UPX�{�Y\_\y��������e&�hX�����V���o輳n�(����Ee)���c�N�M�&����CTϨΊ�{O!rʷ�:�+8��C�Ŝs�)1��q������}�$��g�I�E?��i�R�I�>���Y����.��>�Q�9�4j]��]�iBH���$� _�E��I+F�$�I᱓n�P {���q��7&����;�O� Q\�����y@i}:���(��&�ߵ�G������jv��$���P�}�偕r�O�����yŸ�1|��qO�Yx������,�<�����OC�������8����6���x@4�U�K��7�:�����lMכ��v|��m���z�>z<�$�g��+��6�ZhR����9H��)mN?25]2�]�-��a�P;`���ك}�=_j��������p�C��Eh/]�xw5A$ο2��sC�$+Jpv�{�o艴A| �58�)"�}O�#�[���r<��"��	]:���G�iH�� ��k��[$���2�������SXã� P���x��̧�o�E�E[�8��.�p{�bY����ƞ���֤�d����u�'F���-.�N�Y~C�e���騟���m�9��-�h������4DN�.Ϟ�����P��|��l��%Wt��Ә��t����󰣌iTv�`�ܱ�!Ȼf��N���ߡ�B���mg�tƙh���;]�H��Tfg{�tm�@��c�io^ԃI���73,�B�mTs����Z>����zu���wo��a)Z@�5���������s.������:��׿���vT��д�_??�h�H�j��.�%�ڣ��6���m����z9JRն�HD4�8�b��Wu�lo6�N�)�/��7�*1�B]������
DW
<xL��f����B�����a�u��5�x��O�=B~�E>Y:�#��]؂� )�|�\�	b��߳�����~Ta|�!�!��o�_�;��'�*l\7�ABO�=�&=�vI�o�B>b��;����XA�ܯ6�������J�g�²����>�0��~`5ir\�v�=��<��7j����8϶�1H�5VL���c626�I��#��ZF6���ޭ^OnG[ }�y�CY�<]smD�lH;���-��|����S�f�J-��Q�N*��xl����̫~�66���ѫ�w��X��CMFs౒nL�%o�uE�d�������̍2�B�.D��	f��'��WVL�ω۽�o"IS�Gz�g2�J�o]��ts4��l�?\�,��$�G���Jk�d`E'��׉R���/t��[�s��߹'+K8Y�����%�4^#���v�Ϝ���7�:���<�1�����O kҫܷ���o���	S���{4��'�ӁWd�6������ߎ�u޵p�4�:������b�4���kFi�[��1D��GE}�v�C3U	�M� G.R��h/;-B��l�r������+Z�؛.��BmeB}�HF�J`�����oH�3�x�G**�v���F���/��_}«�%lM�8^�5�#u���p���Jc�0�G��c%��|��;�F�7�,�b��C_�<��)1�7p�o�a�{e��k�D���슽�?�v%HQ�<:X ��Ɩd؞��kZ4'��{��nʄB;��vgD���ܫ�?�T7Og�n���?����z���l������47a�O��!q�0�n��xIFo_�q�uOag+�vMâ���0�(�ϑ�n%��W���p��������#+�Xd!v�^N۞�2N5�dX:v��]�<i1h���:]�4A�SU�'��*
Zŏk���<�~	��\Ğ+�[���82^};W��>h�B�}��y�Rf�4&�q~kX�]>�"�n}P���<\3�n�]����0_�����g>[���e���_������w���a���=o߳OTvo�ߏ^��}�^}AS2��Z	�ie�|৫�	*V��-]y��$���}���H7QR��9�y1�4D������������o�>kv�ӳD��{U9�X#r܍�T�m""�ޮ|�V�A팏�/fх�-���K�sqIģ�
rԍ�6��Z�������em+F�Ѷ����b�����oeh��i�l ���O��6�f�	�g���[��fY<DJI�`����\�S?fP3{w"3�-���il�'��8`��g�ۊ�9$���`�8�W�+��+�h��X-�Mⶌ�:�)� �j��Cϰ����� ��ۇ�KR��Q6�e�Ԑ����#ؑ>��1U�^h�4��_O@����S�_����Gv�zP�������de�Z�%�` �K�zw����gl��+�%��D���O	�\:����#�쪲|b�_q�y���Z&��Pv%�l	���_�x��G���ϵ+<���c(#t`#th�Pka��O���Ŵ!p��f��9�bL����:O����b!���f���vl��mj0B��3;i����YN��9!�Kx�K.�-P�%��1��Z?��\�������rjw:�8�'�?�`񪼳�(�"�j�a�lZ��ɗ4�"G�38`n�J<|#�=��-���xD��)ȾY�5��Y�s�����d�RI��xDCIQ��Y+��>�ƭwq�d���o����(5�]	��2ҁ�⺑oy�Ȭ<��,�/.|�^o�i��1%��%��_?:�c�dnZ����]��1��n?�	�>
=ǎ�x��mOs}��_�ZP��U��8�Z��査���49����/�eğ]sŕ�f]K���̴z����F~�п}��!`�m��O��C��뜛5��u-�������(VE]�f�&d�s�Fk������Լ	"�o���L�rU	1O�Ț���,��"���a���A�˦�~=�X����[pߤ�d�Tѽ$i�¨[DR�f`+����l�ON6G�2Y����Q�U��׽
�\��#��L�$*��v@������+�Q}>N�B�p1�	6�<���r��� \�_��}�3��������~_���Im�P7n��52�&ƕV	ڿ��g��4��.p�����
�S~8��72�n���e)���s��Y֙wk���t�0�s� ���=��MLO?���SEJ�su�\����q���� �B$�]��^�XB�l����YG�b���(9��EEX�N�������ai���ܒg�K��G ��tq�#���6T�*�4>��/ޭ��X�`h�iD�;[6V�q�G<�?1D�r��?'Ύ飘����?����W��G�����C��޻+�LT�`h$��Y� k��>�B]�Ӂ��OV���d�=��13��w�Me!�$|�K�����]���D��$�XQ��ɐ�i.�`��`������z-�y�k)��ۊ�O�5���/�1>]�ū��~��V�����آp�Jc:򎹍ѩ�c�Q���S�C�p��|��!��n�qW��yVnl��3�Y�+]u䓔�9����_��1���w,�D}����鴵��6}�s%C%�l�;�b�p�m�&�+fB/ej��ME��.D^dG��4Gg��c�r�I��'j�_m6Rܕ�lѻXE`F�7꤬bٹ��z~�k�k�ަ��B�~0�F�P�Ģ[��' >b�8�%���+��d��7Q����S����t�eu(j�W�*��%EU�\�l3��}��xWs���'9�r1rm�����>��F9p#֩>o���˗B��r��}��E��i��GT���R@bP=pS*���_�ں�^��Џ�����r��-�V�צ�g-�0��S��$�6�H/�d���k���֧�z���m���3�f���ڱh�[�j�r�u�]�2�P�S~�HC��@`�����-ˑ���{��w}��I�V?�˹w3C��/���f���.��(Τ��v��_�.�^]�D�g�6mY{Kg�$> �J�8T(��cJ��bڱ�/.S�p��.�tC�*�쾓F�08�۷]E.��;��ꐏ
d����V��%�T~��c�ȨM����M�L�H�ϐQ_r�f�D�O�$�|��Rv˕%,'یF+[�/�d.�)�(��b)0	�/1�k�w�F��G�;b���N.�|�z��6�vh߈�����=G~�H[`l�G�.� Ҽ�\Q�5�,�X�Oj6�]rр�n�v��y����Lӊ<��d{B�/v�����ü�������^��%-���LP��ϋ\�+���f�����j��I�8CE�j��2I~@�޵6������'��3��^��	8؋��P1�N����l�6���jKߔ�Eh��^w��d����ٝ����h��*~�4�~o&j��A*��R�(p���3RI6_"y0�	{a�(�p�V�p(j$��C���=_ŝ�g�쪺/���<y�Zgk�9AvU��;���n
�i��Ӭ� �X�?F	�N4���V�P�KE�t>�W��H�M򬚱G�>��:p�g����5]o�����.L�[�R�S���Ѧ�x�	�a�Q<��ӭ���$�)�/�9ɽ�1��Y�����b�$�=Vd���W�#`pD��&��^�5�[�{�0�����f�Td�|^*�ǒN?�df����9II'��iR+�������?Z���&�٦cjJ��N��Qt�>��?�h(S?T���^b�Ƈ�[�Y��č��+�����vJ��?��y�Vg�Y�>'}M�Y������u2���2M�a��}�(eÏs��+�/Mg��>/��N��єhGU���5�G)Îi��mꄝCxa �G��E5�_*�g��W��dN"���@E���C����B�?�t:��B�P*V��g�o2�������b<�t~@@�g�M>�E�r:�&�>O�`!m�����Jv�2�� �D�N4�m,}H��$/I��3
��J�d?��d����'\dEк��h{̱�i�u�P��U�<"S�8D����@B�9�BPh�T�6"�X)dcT{���*ٗ�6�z1�ѱ���1��9 �{�r��C��f���f�tS�)�$�Z��r�����~��Rxsj2�n��G�����N�ױ�����ž����N��r�
Vj) b������',��`+��L�J�/~>����Q��M#nyF2��d��\�D���G��@�W�z���@��o������;m̷9ly��Bҧ���� v��}nu,�$�����*t���T�|e�~1j�x4Z��yT/�jP�8n����h_�d�Zeڞ}�������<�e��]�r���WM�?-���M���o�%Bc�ӳd��A��42���5+[�?�7n,%�'�߰xx�v�c��x���^Y��F���ȹ��#��[�)նvc����/_0��P�˯�J/|��%Kf��$�r�g�w �"�(����6�y&�$f���qy����xິ�*��7��F�*F��E�k�O��3����
�<8�B`͉m겫�h�D�Wc�ɳ�)�9�r��t
�J�e]�~�Uze����#mqv��u��\�N.2���4j)����:���a�-<sn����&��4GF�LR`�V��`���J^�x��Vv<7���/�u'|*�׿�����.�����?X1�����6���[���N�j���KG���p��4�_԰.3S�c�>�X;R�w�vLǼ��2n������ʘ5���麿�������S��ˊ�����t�zs���{8f�n�6�J��-����z��]|��+'W��T���L��a
k�=�~�7We�c�R�/3�>�`��ڏ��u��G<wӯ�m�E���G�g��_�7�w�3� �M��݂��)
�n�[҅O���;�9�і�=�c��"x��x-{'��*���*�H9L��RnA�i��,
�҂��oJ���M�RD�G>&�hk��$-��ԡ��
wG�2�u�����i�z��D����B&ǲ�a��~�_����T�Ӊ����w]ق�
�����{�C����nF�d���c<%�d�������u�^��/M�T����?�,}P,�X��/��,͂<93�5�a�g�阽�ȶ�8���|�8�}��Mc�\֓rq��׵D�����A2o����=d3.�=&}�6t�s5��ֵr��'B�w���Uޫ �e�MM�a7�����[�TV��ٔ?�V�b;�C-�t3���N8��UYT�3s��_����ܼK`Ԋ�}7e��W���ttw��'�-Iz5~C�H��Sv}.Yԩ�;��Ɠ��d8��qM3E
/1�����ng�>��eL�������@=�����^����_���~�0f,�'W���~�|FPU���S�� ���y��=*_b܇����	�MC�v��ڭPz����o4�e��E��K�Y<Q����yI�n���Us��	��]h��n��'<����5��#�P��O�b
Ѝ�,����݁ �X��U�QQ���}~4�4鎰�,Uر��G
G�,�zK����ux���� Y������J/{�����;zU��N@����E��^N��J �N��c��j�	����GJ���Yã�5W2�D�����Uվ<fc~0�����]��k8����|�Ft��f��zʒ�
\g0�n<ҽ��I�NNL������L_��0�����q˃�$@ۿi�*Md�XA���9�kr�}mGF�Ę�	�B�7�z���X�F����t�W�n���J��ѽG�)�cN�['H\�:�YX^��:m�0-|���r�U�5oT�=��a11߁���u9����m���K��%>�X˛��~��7��L�Y;DgX�[�Ba71"4uh6�&����HE.��w}�k���+���������������}�8;���o����x-}v�6�ΐ���x��[�|�F�꤁�xj�.�1�:z�9�y�K��Y�'��=q�{�����ߦ���3���3�6<�x�-|����n�	'�G; �-  @ IDAT�����8�ýa�.���_ҿ�����wn1S���/���_�:�C�dP�?fey:�]Zߚ�Q��}1�;�g�1�ih�:3q��{��u/E�Ц`b�;-1�`�&a��mZ%����	4O�SY�8ٍ�R�(�d_�4dY,�IOG�#��={&#��m��m������hKW���81�8���3�G1ӌE���M���
�w]֗�$�O!Xg>
�:;�"_aLp��q���5SZ_��_�7�F�0�o0�:<k�fq��=��)H�g�#j�aN����]��i���#*
9Q��H*�nْ��gYɶ�����t�����<<�l�Ӳ���}�q�k&����~�j�{k������1���I]�SS�#�(t
K�K�E�EY1�Qڅ���	%�r���q�:��xth��%�u֕B���zBL%	�k�֓'ͨsBh�e�\�3=�s�!�q���S�Wq�v�j�@I3^ӊo� �J�'�i~��p��IKa����� �Q���7(�Vf>��/������+�?~����焦{qZ��D��/Mݓ��f�}���q��1��*����
{�$~^�Ñ�*���R�v��ff����\�Qw�ғ�L�%�f�։��-N�RNXxm�?5³ܸy���1���7�tA3�R���{4ǳ_J'-���g:�T%ei�Չ���S'�����W_}��?+���`�]��#���4��b��ӷn�P���ĩ&��R�i�>�����x�:�B(ݽ S����e;��Kk��<�kP�+�T���
4]�hϱʬ�]�x%�=,���g�G쭹�A7�+{�!a����*h�ҪǸ�o��~��������Lo��e�U2y�8p�T���ZP݆�q��3f�Sˎ/�N*�fshT�#cU�cb���|D��@Q�둦��G똃�\6(�<��k*C¶*��+)*Ԁ�O��S�4^��N�x���#�4����F?�@��zt��QN�����3����K��oӚ��>��_��0��s�����W���黗J�:��[	월	�~��ǘ�q��m����ʏd(�E�Bk~QWQmbc �?o߼E�=���&=��W�'h�,�,�VF�T����ID��k䈲���g:��(�*��3�~-�#��㘺���r!�Q����w뱎2����xjﱡK�_��P{�<���n�� �ŀmy�L2�.��	�D�(��֏N�qa�i�y�'g�l��t4333������{�J����d0C�3��qٹU��{]űې���k�ӏ+ h��aO���]0f=�ј���Q7=�q��p�O���n��9�Vw��v�W>����mi�w���Oi�&*�P��i3X>�fIF��V_��j��4��^e�6��/�Ӓ�Y�8p�Y��j��E���u�Ṯ�p��2l����������NI���v��`��W��q�r��ر�u���o�N�3h�j�5�F�-7k��V�8֖��1����� ���o?2���y+��7خ�O�%Z�	llgo?.�~�C̖.?]D�����Ux�L�r��j�����B9��"�ec/���t����)�y�����'�~cR�f�AVk�1�~���`k:���=j�T�cD`�sԇ�F8ɛ���A�@lm~נ�8ۯ+0�#<�5s �vcE|�����&��a�	�e���T0�B�^=e�̀�|�.�:x���TԖJƈszz&���e���J�wQ��ڙ.���\�^ƕ~�*}V\$~]5��k��n! xf�p��<z�������+^�� �/>b��g_A�G�Yk~����
y�п��+���~#E�w�Ar�y,���?��� �8
�k|Ϡ�S��GVY�Y���o�]C�����3X�i�㠝N�!��vCd��f�f.�%� X�\�R�ߤ}1V6_�fn�Xk�t�>�	� ���Bv.�Wm7�� �i��|��ySr��_O�r �`�Q�U�[�J��ј�=���_�~��2�L�?��|Gۿ�՗Ж�_#`����� ��'	a��6t as?+���h��Y��oО����n��*[�7����Kބ/7T���8�	�s�~x�N�zY"��@<3��7 ��Ky�O��5��^ĵ�m�=+h����2����aN�0�j�-�ET����VH�qS>���݈g_AD��^a#���^����哏U������e����͹S��(��"��o��~ѯ\kƥr�
�J��^8H��qݮ�	�P!^�[�Y�0����������>Zd�9FПxzVY��CWqF����{q�1���QO�Z��X"".���D��d��#L��W^?���� �Q������Ϯ?��p���L}�7�s�:��zw����"f?7D���_�����rEL��7�$Œ2��YE��H�8��~���p�ϡ�
��c�A�)���N�Y㛔Q��P�2���Y��k��E�y����z}�����ym���
��#�I��g˨�Y
���c�9�`No[o.����+��~��V>�3?�M+Ӊ[��_'^�m�u≓mOW���?dd]��������\𝧖}���<u"la�G�T�j�k�����Qh$�����:�T�z��C|����̘�T�G;�δC�$f����$joY�x�a�{¨pꬂ��I�e�>s���W�`O�F�ǌ��k��׿���bsM��,�*���6Ͽֳe���g�1j�D�젩�����ƻ����ǌ�>De#�y�&��_#D~Z.�Q�%��=1F�m�!VAw�zJ|W�s��u�@���Y<��	�+L1h4�v�^1,��?�O~ǟ��نX�nZӀ,~nJ_q�9K"9��=�g���m�����y����=�Sc;A;<���Q�:So�Ai����tnr�� ��M��0/��6a���^�����]�֑B�'�A|7���$N�Y^�+ݶF혩1�*����C�Fx���_N��x�̜>��3�I�D�`�{Ʀ�uf��Z��ɻa����@�hb���S�#��;����{8�+8J��/�W�h~��#��`�=�L���<�Qs�#J�x!�8߶�`�U@7ZC���Wږ}U��mz�kư���Ĉ���8[F۫|�
���y����ô���c�B�ߕ
�;�c�g_',�Ȱ�'k��KSӧ_�W�>�g�s�a/&�B�����|��;|��@̖��{NƘͼ�)�uf�t�r���c���޺IL�&ؠ�%�>`�Aaf Z�SG�/I$���W�uoH�/���ޠ/W�"�T�\]��#�xlG
lwӹ�{y8������U���[J#~I3q��{>���>öe�9�.�&8xzf:����W���?�D�N<Μ=__)?�����jd|7 ޒ�7n��Dg��<0K����V����J<&�lﳬz�_��W"���kn#�4Ɋ���~X����H�&Ŵ�3L+U�����ީӳ"���\q%��i<��Zy]�0�{6T�����)�h�f����~�~7���ꫫ�^���ܶ����!��޳��,Ɛ�DM_�<��b슅��C&!n޸�F�#L���
�
�)��g��k��!�}��\�;LHipN82�u���B�:GY��i/S�fp��w��Q�ae���Y�(+0�U<݌;I;<�q��e�̭`�Ƥ��徦���>�߶;�]��c�1x.�q"�
,���,_��� �yj�{h���8��1��Y�t>����o��=p��~��k�_�7�����3�6��$N��[\|6�
���s��N(o�i�Wgz��3�E��ۗ��<&�"����6�����_��NZ�媛�jQ~^��\m�����_���BћiV�������|�?��S�?7��a:�3�vg,uY����?	�2�8Pڸ��Oq�Gt�s,[�`�m�.0+p�������?��W�����Y��g���I��"Z���F��w�h@�x���ĩ����|�ɯb�W��ǰ�߇r�*�'}\C�`F��W{�f��OAf�8�H� |`h��{h��0k��9���޳L���0L��6L�|�p��+.pEBmx5)�C�N3L��
��:3�m�@m��gg ~�᨟�h�)I
lG��tp�d�=(���)�o\F �_���ܶ����.�:�:��mm�cIl'��n�\^��a���m�/�_*u�� B��V0V(V�uf���X��#����:v��b�f��5�/�s��a�>�L0�3�T�#�3j�#͢C|j�hi�u�V�~�m�l��OP.�l̓>��/�I?���fO

�wp��¯ʄ
��L>`C�=&K�eW�]�du���Q>T(3���p��wXm�y���/��C�(��Ux&��F�r�	�)����p���G�Z>�?�ar�Pᠸ�e
��A@	r����{;
ţ��Q��O��d-��ߒv���~ї�J;�|"��c*��Oa�z�S��̔�#3����T�z�[�t����~� l����JwW� �E����w�0��l��WU������Ɖ
�B�~,/xd��Bj&��ܪ���&׆]U�t����[!g��b�����Rx���-�sa1����%����:�]��?�3E�G>}��z�����vi���o��@��c�W��'�k(��G.<]�ԋ|��xF�<5Ǳ�G�OP��[7�﾿�F�8�#�J��1�HY��,�v��*p�=�az�e���LM�\�P�t��x��z���W�:�f9�09���k؁�U0W��ce_�.�'U-G�4��=���8��i|M�ȜU�'��y����e#������k�Y|B���> �y����|{��$}������$U ���Q�"�䅛�o�Ͼ���C�ؠL{� �))�+~�e�9
�,V���#�[�`���
�  slvs�
�c|_�+��b��[癃ऺKW�C6/;�o.p�����cZ�PZ���^��۸'Ω mr����;a�u�i��}��CM���0uޭ����{�k�����|�güt������s'�Lg�}���D]'	7��1̲8� }�3��mER�8*�Ʒ_{���RW��D6�.�{&��_��\Y�J�N<����4L��}�m��Y�}�e�-�)�_���Ba��>W����W�����w����#q�L�Q��,��MS+��B����3����~�������*eW�[o���]~�L�i��P t��,��03�Qy�x.����f����e�n^�|��e7�e���)ң�9����;os��qB
��lk�s�}��6��{����:)��X��|�y������T�*+��
�n���ݭ��:�:��y��<� d>鲬��������m��kﻥi��9V#���!T�x u�804ı�-��|[���ǰ��3�ډ����\��3�:?��� ��4�apP�\�}W���3�
�����L]@ig2Ł�$8����S�}nƠ)�Ô���OB�g��v]��`��؜����N�aSu��C�4�-�x)�9s������LcC�j�;��Q��L����a$�4I>�'i���7�� ���0��c�j�8�_i�잃�+)�t����Xe��Q}��*@�=;���L�2�� 7��i���� �����!�ȫ4.���X��1�p
n⤉��a��n<�c9���`۰!����=����G�u�`��Bh	�����6��|(77�e�|��u���v�f�����9�y�)�3�)aX?��e�dSa?g�ܘ��<3��g0��t��q�YG=�.���8�����ml�?����[�R*�]�@AB�ʒGu�����ᘂ�?f�� ���
��A���<�G:]�� ����|�K���:{Q��8`�	f2�����������D�Og�yY��[E�E�qp�=­�x��7��'���p�m���U	�B�0�_��~�9�7�]�.>̦r������Z�yq�/�@��1}�g�u!Ѯ��tb�|��Gl!DͲ�wm�>���3�@.<F���C!�� ��c"5���z�!�s|������,2õ��"����A/��p�ߢ��&������wi���⥐�L�*p�h_���&�d��\=�"�jsH�L�xԵ|5�j�������Ϣ�.�*�ֱR�u�P��!M��ߗ�/_��U�D���E
���{��{X<i˺t?�8F߉l%oo@/��P��K���̫*���z�ѩ��A�o��^���ߗ;��5񧜚.�X�ցx:�a�0M�����&xn�VY��5���U����b};�Ap�w���=�oF��>?�t�p�H����a�հlK���/����4��L�[&�&۠���g/᛿w��Eg��v����Ɛ��u办�H�7�ru�2����v�N��Qt�q�u��x�r�͚�9)uf�t�eNA�n������[+��<�ĩ�z�d@�i����?�p�������"a����A�ݜ��"_�~,܎OXȥ��đ�3|m��w�.'�NE�}ę���8�@�����jopڭ��g#U�Q����Ux�����+G�j��3z����sq��2�۝[�Q8�ӏ{�`�۽v�l����q��B������W�(s�ݼ�ePϽ��3q
�u����c�<�/,x,l~��t�j�N,N���my&�&;���wt�a��h�:���ÀE���]��mG�@\��4:��y�&��'nvƷs܃��`>
P*n�T��9;=����v�p��B���|�Pԣtv`�y��mVz_�x�\�vQ����\���M��Z?���ر:S
�~��Y:XWj�0�?�:���^E��ϟ?_.~�C��W�F\�U8_�YN�u���]�yޓr��rGd~��.��TcY�0�&��1�9��!li�@"�L'�[�I�\�(뇦T��]
�)q��~}���6�������<Vm<Md�=�J�3(���w5D�di�ٜ+�~�N7�Q�O��3��Ǐ0{�%��sff�	�_F�������?F}iN��r�@����U��9'-ͷK������Fć(���_��p�|��s��!�g���¶���y�	STH��7q=~�X� �� ��h�����	���c��)�e��]8]f�&K��!
��u��u,��(����-lۙf�� ���G��ʳ��q#>���U=�>�ͩ'���%���/���{I;qp��y�쥒� [�m����Z�mk�����	�)�+��s���Y�U�z��-����Bݸ��ï~���YSC۽c�����褛f1���˗/.��I���+��o[�q5����Pdnc���q p֓u����U������1��˦s�gX�*֏��?�����jC_�#���h�������<��{��)>���*��a�C�9�GPr�0��_�go�&�������[�/^*��Tڲ��:���x(*v⢀��݋e;�[)�
MĞ
��T2�u��)�|垢8���VX�/�^^�~k��Xa�{A�r:�)]��9��2�7|�,�8ۥ��)J�0}�}��+�>�!k�D��J���W�u��3I51��?���&�F��l�܂�9�}�э�u���,�m�{�����Ƒ����:V���cz�gz��2�����0��p2�M+��3��3<��x�K����c��S��u���5������M�0 ��7�5m����iQۨe��p�cq��7�)Wi����TE�����4��8���e��my��%��_��_�����3�ڹ׆ee�!���m�V��-��������Ͱ\|.-����s�'�0 �>u��a��l�|��8+ze��9qɀ<�Y�U�-G�뽷\/��x�tb�~�{����8w>:�{���o�������H9yb��j6���|�3A�H�'F]�e������j�ƌ%�N'!�� ���ϟ3���C�P1�6ݙ�+W�!\�N(Y>�k��{fx�2n���~��c7��'PG�}**�S�OŬ�3t�j\Gxq��GaP��N-�]v��5�є�˲*��1ic�v��!:�S��<v���C�SU����/1��{l&se`~P`�q�`� ����1�u��rT%g��� �'M-2�|����K�qz���˛�=ʌ��|θ��3������?�r`�:9wg���p��{i�/��8�QeIS,�Ǘ�+�e]{ϺM����g\��@c���@
�~$�(f�;]r��4�Y�ȻR']������7y,2�w��<�͘q@��gߌ�Q2��4�ߛl���VwV��S1��o��Ϳ~�:�w"��t��iu�\�� �7-�-s�?^�kal_�9x�P���j�~�~��������J;crV�zi�Ү�D�1�۴7��8*T��A��1N5�r��������e/�i�=��*F{Y ��
�&�/?�"Lz�O��2�d�
6�����k���}�q�Iځ<< �✨�`�2�z�����hw*��k�E:�b|G�|��Y|ۣ��7�;7�^E`8t�I�#|��7�-����ϰÏS��1�(�*���໼t_�'7iG��p�I�H��e�G����lφ`�������(����ц���ߠ�J��$|{�mz�����B>@�e31B�q��~x�n�]E��8��j��ɧ7���~���K���
�<k?����[�6(*�ڛO����2�|�{�2�L���6�q�,
����ٳa�o݈���_|�M�4iU��ž@�Y�ޥ����g������op��D��/h���
�	��`����4����M����V1�%�S���6��~C�>6���S�'��x�/o����z����S���d��pY�����ӿ�>ҋ��5a��Y&��?�&t��v�n��)~~�}	������ܛ����?����-B.qs���(�s��X�!�ʼN�ʺg�1�̙iV��p�.�ԩ{[T��O'm=.��2�
��t�k���¶a���u�Ig٥C�U���pV�`&L��0���,�$���'��I?/߽t�m�n�*����8o����Ё��l�?��|-aR�E�����\��~@Z$�,������
auU^�O;�N��;���s�OR(�2����|��o�V��?��|�a��XY�(+�� ��y�܂�g���(���'�!�g����[�P &���f�i�YO�8D|�:d�e�&�f2ګ���a�y��������3n��`v�؆�G�Zg����,�}/�s���hy8�2����C�ej�d����D���0�p{��)���@��O�8V�}��������e���0��n`�QΠ�D)t���؞�WY�6Oa[O���9��t�s�����1~t��]O��������8B��I�u����b��1N�9U��NEپ��kNA�'P��&N֝W��0�3�E1V��}�������٧���5�`m����SGV�����Ry�̪K���Ӷb'|�IUPM��]g��r���Y�t�?|����X��VC��u��[�QN�D���fEQVT"���e�U$�2ˣ��&:�b��<I���36?b6C<Р󮃐����I~��v}/��0m��	wC�F
�**6�S�W�����Q{fsȎ��	'�9By�EM��ʵ+WXqzX�#pjg�`;�9���c�(W�<ޏ	R�P��^�&�X�4g��=/���_`&V�qgu��b�3��nµ^�ێ~4ᔘ�q�Ʊ�7�V�Cο�i�Ҡm��h�c\��䐴���͖�� ?�{����[���*���N������O=����_G��!����@�L�c��V�B
3�����/�(y
H0�����B14��~��oJ�`��_�.+48ΉW�����+y�}6�ax���2�1�!h;�����F�v�x</��ʅ���|\����v��u�R�#imy5y2,馟.�p �t���%­[�A�i~��Mc�/�>�#�f\�~�4t;�����BQ;���i�_5�mOr�a�	O��`������x�6)M��U��Y>&�ʼ��'i#�P?�(:�]�&'J��ҕ+������+����j��D���������2k�L�����se��QO\���7Ln�Q��2��1�Lx�n�u��6i��5�Ϟ���e�����M&u>��KVU�P0��ǿ��y�S�)�����`2g�U3t�X�������J��o2��di�6�ާq��� �fS��$��=�cH��#�N�X�q��β��1���v1�ʉ��2f�����O��H3L�p�;�E|�x��)E��a��)O{��X���;��nڼ�[($�OX�pE����3�p�$�kF^�g��1�-�a-�g�d=7��c�P��G�x錛y��|�?�I�<!���%����*�	'v~���_z��va�04�R�W�p���~υ\�@hk㱢j�ꤡ��N.��EY�����ܝYvUw����f�Fb2.e�\����^����U�ݫ�M���l		�R9)�!�����~q���T�N�w�9����3Ok��z�Ҕ�/���F�K����w~�^mKPN��şf��������7���q��o�A�ӡ0�i��?ef�/�����£L�d�ѣ�驭߂��&���?�=�O��?�!S����Ae�;-�������@3�� �(��Q[
����������2�g%�ǵ��{�å�q�|���'�,��KF��Stv�R��
G�Z;{9��q,�jaf�Z�*�2�oqU&��]���|g�������7��Q�gҘ˨IFʬ������7_�}Fߍ:����W���mx��o~��Ub�B�[��#��������6o��Fe�[�s�j*�^�����rF�����s���������fm����G)��?�ܻ�����4���3:�p{)�EۅJ�Dȇ���;&��￟�\�JM��uN3k
���^�����L�7�������k�Z]ih$/�s��R.h4k�XlT� �8M��vl�-�^4�\w)����I?�������M��.FgO����9����ߏC�=�g���n��N��]a�ɱiT��c)�_�..�q�lv�87��3z�����tÌOF�"+<�[��%�t(�E�pF�96�4$�X��
ى8�<,�.�Cד�v��s�T�`&�U�蠵���R?��?F�7��7�.שv5jW��Y��:mʚkz�'�Rﾹћw|��������E�N�S�����,���,��9Krn�gS�i�4Q%h$w1z'��4K6�}b�\�Ddy��W߬FBR��q�Ur���ŧt{���\~#����\֝��?�0�c9�t���;���:���͌6�R����_i �q:Ɯ��={�=zF��C^Ҩ$?���䏟��'�������}7������Ϳ��?K'�e�̈́��Ϟ��^�B�����9[�{6D��K9����'�	]U_ՇY�%�.��n�����:�Ḻ����t�!�R�$�CӅ��+��~��o���'�90*���S&]�8z}&�b[B�u��'nfpO:MZ��f��|����=a~+�W$����m �_�R$�b�;���9�Ѹ�s�����l?����;Y�u%��^eYo}r3z���tk�{��3rAw��4�SP�r�1�:�sI�'��ä;MҰf>
�M�K�OY�t(��(��=W�S��=J��������S�~���/<���r���;�$
ԀB��Z�_��[���}�:ZQ`���<���7ұ�ޢ�K�>�����`*��yҪ<���t�=p�&�ox����+'|�u`�M�6�	�����^��W�pMg���t��<���O:e`����H�X�y��,	�����L���s �~�N��>�#3z=ʑ�u�Hfٜl��u/�w���\��M+�03���I�&�_~pm����6��/�ϲ��+|���ߣ�2|1���N����I���sx}KH�<��l*�6k$L̺6%[�	�4�B2������O��'���ԕi���B5���CG�c	�Bߺ�{�4�|�w�������:��m)E�IL�#���w<8}ϣ /|��*��g�z��+�R�85�T:���9p���Y����9R�0��\.�y�չ�\Gg�9�t�|��i���_뢗	}�2�N�'Cn�S�d�P%l���_ys���4zގ܏3[��͇���$7Ҧe���������훛��?ɕ�9r3�����3t�%?�������*�z��b�t����}���o�.���4�2�j��{����Z�d$�V>8S	m���_������w���K��b�❌���(�Y�#��+ل��_�1n��|��̲ w.d��?��h������oi��X�I
.���|ms�g߭�Q�b_�z`i{-�5ꮾ���Y�'_͆T�@2ä

���Cc�4��K�/vǎ4��K�4&�fZ�}��m���p
�эo��v�E/_�jFy3���(�O������ϗrg�w����뎝j��:�tL�S�H�Y�<iraIG4l�����h^8��ɯ�LM���4+���I��ɽ�����op%��עðZ4^��+=���f���mz!Y���������܇�MȌChڐ�h�.��/^���'�,y8�Xq�I�^�TN#u�����P���oo��|e�q6�j����;�rJWl���-?�Iĸ�Y���F��5�KeWG��.��Q:�K��s��)�h:���e		��)/�g���_]������_�����_�W�x��cٛu�Ƶth�e6�F�9��CF���%/��֨���P��ś����r᳔ ����bY�?�K>�%yk�
\�𷧈]���4
^�Fl3O��QЙm�������3��n5�ѩ�KpH+�����`���X"��I��9q�-�h�^�o�����k9�+�&<���.��,��UfI�|�k)/�(Kdz��>�o������7��4��Ϭ��������iʖ4x3;w.�Kt��/���2�nh�=y�+ݍP�16W����u��&#G���C\h5\�ٯx��n�NG3˄<�d�{����gHn�;���~����4��� |�Z�%o�g��]V���,w�6Kj��?��_�,����G������<��|�Б��N�������,�Ǜ�����s��{��8׃��z�D?t���>vݻM�AT��ώ�x���/���p9�+2�%�pt�*�,i���Ћ�J�:�L���?�]���>3��9�78��������K�h.e��hI�t�73Ș���9�W�(���l�r�~-���|:�aFZ�hXzJ���M��$��΍������]�iWIG���H���-X k@o�<O���|�C�S�<ɴ7�ѡ��j�?:����,�{e}�W�	���t�����ѽ_�M��\ܨ�#�ذ_8ti㚥>o&.�M�:�d�g7|]L�|?K��h��&3�'֌%�r�ߺN����~y:��n�g�(w��X˰8�UU���7s������t�_������\�� 7�5y�_�ǂ��gq9�e���(��eFkn޼��ۿ��l��/5����	�Y�s0��<k��ZX�C����� >>�;J�d�6�O��o��S)�\s�Fp��+�����F�Wh��B���,���e8���������1���b�{�'��=��p�9�5m��96/�o3:�z�id#�p�p1�r�s��e���ܓӌ�0��;�df��.�Y��/�щ�T��_�w|��l�2���[_ΨGn����_��'Y6���;��A��O'O�����3�?��[i4�Q�%����8,��
o�)ֳ�W�����J�x�,���[xU`���_�a�WA\�[Î����TJF�����׿�vF���4;ݼ��_d�r6ܥu���qN�I�u-�qi?���揿���o����1H3
�V#�i�(�ko�}��4�l�>���W����>7�H��F�4F]���/���ψɫ�+�'���3�����/ܦ����ZdL�Wi�A�I�;N�
n������_�+�f�O��z乑e����|���r�����~i�a���K�^�>�55�T�x����~,�4�|�{�����qF�3�,����/3����'�5�RVhL}�MvfRl�SIܽs�f��|���pLŢqԣ� �'�O�I����&�w��2�+}<`��'�T*}���p5�1��/߯�
�����̑N���G�J����]�j�_��>��E3�R�Նx���w?h��X�k;IWK��~����ַ�8��FJ��N�����ok_�^�"e|��ކ6�_���W�y�F�F'�ǥ�ˠ�8��8q�u���-�f��t�kd����t��c�¥\�|w����88����Y�sy?ix���4���J���y8���Cs'7��r�O7d[�|��q����ed��x��������Ʊ�͋�}���6�Er�����:A)����e�Gy�'�t����T����K5�;��,���GK�H;�R�����$���o�{�[x���r�{Y%���׿�zJy�f���Q�S���N�R�c��u�N�j�<��[;a�N&F���^�@䩃�}K�r|/��z˽4/�A�>���^�h�NNDět����~�v�$�с�:YliO�F�������1�|ay�Vӡ�GΤ.�������4����Nr�<H�
�p�#��23���?;1NY;�[�8��8n���P��]�n��1��e?��Izy�X�&�%��<���K^�@leHy'����L~}���Kcy�1�O�qi[�|tɁGҜ����qp.��}:ǹ���".�V?Ձ6�0so����Xn�Nfu�V�[������s.m0�|-uo��}!{W-C�r�@ˁ�K�ҁ��uI�ĂqߦKT����_�e�pr+��g3M�����Ї�;�Iх
!�-$�8=�޿�bP)�R� ��(�����4�G��__H�|�6����b�F�Gv�.��%Y�FyW<qǕ�qI��]��9|����\�����&�ޛ&k� ����;η�/^Ҙ�k)���J6l�������S�eܿ��a��3j��G�Y��d&A���/f�dpZ{)�<#�on
��<��.�h/)���N���ƍkY�|#K_vcKY�u��6������4@"c
��Ә{�+_ɚ�2ڶ�1_�6��]���̝�O��%��Kc�1�5ʶ����`Q
ȼ�\ʲ9����^�o7��_�H��H��+_�H���G�� ���չ�tȅ��<�r;Ӥ�r���|���W7�x�+�w�a�~�v���l��ӡ��@�sq�Y	i�bW�[�3�鷲D@A���"�T�V�T%S7��M�=
�k'�N�`X/�UZg��⤃:q��Хo7�*�J��&=���?�^�_�މ����=�ޝ�ů4A�r��_�l3�-��~=h��M��><�|�}acyR�'d	�%EN�y1��k^N╯�Z�F��Q~��q)��GY��Mة(2^R��̓/�8v��'����Q+}'�4:�7y�yN##eמQ��;����o�3�ԭl��8�(���2�7ߪ��k�2�4���_x�J�^��42����ݒ���ek���[;t�rF�:��6� #�pl>��4ˈ�%#��[{.�2�˖[g�`w���t��!�U�/�ϧ�4��/�k�v�V����0N���kY@���0��of�?3g�?��{d�p�=���M>#��J�A=4v�u���_t�5m��AF>u����,��K��y7e�k�����_(U�Z�RzK��կ}c�0�Ƚ,��A��KYnƹ�x2�CV� @㿓>��,}��\ҁ�i��5]�e N��D#��^���rpNY�{?G�
s����uH�x\�2�7��W����s7���>[ggu(\-S�^r��{�pxb�;��ntk���i|x.����r�W6��,i/x�{�K+m9auz����w´��
�A���_�I=��NSN��F���S�W��=l�?�uj`e�4ēO�xH����+ـ���_�8����"w�4�/t�<�P��k���ܭ�����|P����-���:m�粏�����Y�D�(��8?��%9��L  @ IDAT�`�'�g2�Wz˷�$�{h]g�����c҇��n�ƶ�oq�]��?��}l�?nt�~0�C�>�<���ϥ�z6ˊ�:=�׼�%k��}�!;f?��g2��ޥ/�+����b�����>nS�Uf�d�W�Ĕj�ݚؿ��M�tu �u��>�m���~���G^�JD��7.l,�#��M�	N�*pc�6/�f��M^i Y�i��t7�(8
�C�)�Ç��9��[�W>�_Z�� ��٨Բ���/�q`+�b|p�%m�	x�{���K���_�r��T���y��+�Y��t7>>�ȋK�� gM�f�%�x
��@,��=ߌ�Ɇ��:x�p�
_��Z�p>C�A�H�{?���4ip���K���z��񻙵�����z�`󕷾����e���H��1��ЌLË_�\�5LX(���u��M�tcY�vS�82�� ���K�����m�qF���rʒA�9�2��cF������KV{yn\�U6���,K�ό����5"&}c�ɗ{]��s>���}_����Ͽ��ʗ*>88�q��|���C>��
S˭T��ˡ���U-�"���n� N:�j+/,a���<�|����?������ʜڟ�%x��˻x�� \*����T6h�;�&?0�K���~�΂���f�����Ne۳��~xСvoK���;M��$;����E�6��uaa�q�_�p�_�	~<��$U���
�fT.����#�p�����N7�fc�SŎ�ٕu$Eѵ7
�ѕ��}��?�w�P��6��Y^���ͅ'4�bY�n��|N^u����7��]z�W�Ý�t1e�q*d�TN�S.���'I3r�_v5�� 72�adt�=����p�l���I5���_x)�9Jt��G��]�F?�+8~�����f�0����6�{!��5�4~m�>���;9T�W�N�;��K����R����<���ޮ���g�ٞ9�^�|&s)�y�8x +���0�I<����r:��U>�wtnضx���|�sz�nf���Axv� ���M=Ħ�y���R����?Qj�鿱Y�O���z7��^����;{�~���끯�K�M�����p]KY�ds�n���#�苝�;KS8�}��R��)�";~��;Ķ�PM<��O2bv�c|��>K~��'�{t�ޣ'��w�N�b ���
/e/����
׳?�s�E2rͶ�&�ͅ)����ËC3�H�9�]?NnGf|���ն����n�eM�ai$��iJ�ҫZ�p�]O�����`�F�Ȋiz1e�����O�W��#�pV^H��,��J�Q��9���!�M酉�ݔ�X }ʟ:����9l��j��)��Yr�+�f�)?��r�.h)
A�"=��W�2����ƻ�1����r6���9	�՟�;�%?N�	ѓ2ǘb����(�sʊM�Ge�z�r�����n6Z=H� 
:��Ȣ���
ٞ�{��/��>e�Q��KJ~:'aD���-�4U�%.p���2L��M�o�/�̹�M�-4Z*>�4���]Ѩ����b��pƾˈDP��;Yo� =�s�f	}��B�I5�f�3Y�J���^_�W��0,݇�H��.�u�����ߵ��v)�3Z���˛���L�?=���9�"��;��9Kj��^�����6���HI��`R>r��P(�Mg�>��.ƞ��[}{�����-�l��s�7��_Ҍ���inյa���_�;>��b�$�B�x=~���s�<��O��E۞���c	-���;<���aGҕ��^�7>�Y�+��6���f?#���+رq߹�f<�#A	��K�"֜eh���/�#|��ǅ4x��?4״vҢ��]�_Ȉ�%w?d�xp��F�̚���p�-��<���~cp-cu��R}����͝��턥���e�\L�(�;)X/���S�N��(������-��ɧ�3��o�ՓJq�}/+y�3k��_�ʍΊF�>|HG�W��WK]���I���c�um?[ip&�t:`����9�c]&��h]���s��%mf��(�K�~�5S�][E�R������\�g�}�M�mx.w�w�:�7�}�G|�p8�?q�jhW�ײ����W�e��t��]u_h�Ђwx�N`¹��^ˍ6�g4�O�i�����s]�j���t�SUi����:FN�c$��螌�	�7���J���繓E���;<:n%7�W8R.�-K�F�x���߅t���Ɂ�C�Q��|g��z��-⌾���ٷ�)�z��o�sVV���7Oɚ����-�ȏ<;˒��ʹ�љ��4�l>�:j�r�,[B˷:`��y��ٴ����\F37<�-�ՑǏsq�+���Y�W
v�W�iʐ��at �~��%��FK��H_C~<r�=������P��}�ɩɻ����.�WfMþf;����	.t�mqƏC��/�$/�,�O�.'�?c~��������mh{�����f��$���f�e����/�f���Χ�~�qx���K㥗K�=A\:�囝����+CNGk���y���~�����{5K�3Li;P�)���G'��YCx	��t
��}�K��υX�'Z��j����2���F��T(��9�H�n�?^
�t!�Os�LF��u�/<�Rc;ʺw�uX���[!�G�?z����p�6��l�����1�gZ�T_�^O��ʩh/
�x2���#�zĕ&E�k�����w#����������ۙ1�1��g�+�*sw���̩{�ҁ����oG��tƛL������U� 8���+����H4�e���tJӦ��n*�'�6���3�x��/qY��J���d��I:IG3
d0Z�EqRMmz
jzl�K�.L�O9'=�"3uE�a~R'�8ictJ��)���/�ע	f�n�q����9y73f>�f���Ǚʿ����>��u���J>�?1+�Y�t��d��"���!�=�F��c��.:�ӀL�������u/���n`��~ů�4���C��hLoa�!�.�qӡ�/�lvt�,}�$�P�I�t�a� ��q֪Kypl_|3I������\�g�.����!c�T|Kq�0b�Ң'�NQ�_�q���mp���&]8�'����{�'Tֿ�XE�~�7z��	��o=��K㍫�?f��Ѷ�t��HF��Β���k8�=��w�����Ņ04������8���`,[�4�p!�����H'��K�����br�#>8t�gs��^��t����8<���3�[I�J��ȍ�0r����9�Ź�#�����"rt;���3���u�Ò~��-���q��~MZБ4���A6zFV3l�O��N©#��g:�Ч�s���t��L眮�20 w����#�wp�At=�T��=���_�$p�r�F{��h���ɍ�]��`���~��>2;��x�7v}��?����~|��� n��w�ܤ�_����o�t�)�.9I�r��C��4J������	>_��������(yn���_����pE����N|r���d�[C;:$σOj�ݠ^g�� �U��4y�/�:|����[��ٌV�������y|�	Y�K�`��-4�0��%�y��Ο��L~�[�
o�G�gɪ���#�6����"�����"��N�����w��^+m{�&�H{��_�2�)~���7�U+St�Ǎ���Yύ����@gk�~��?���k���h���79p�\���la$���z{������M�>k��X�֑���M��t�\�r�}
S�^5N������2�I6O�M3Z?���M���0#��%Q�����?��`@C�p��i1~Ʈ�R�q6���Q.z�(��$��O�:e���Ct3g�[�nφiLg,盧��Sn�>��;��s�Om�J!� �����,'�|�e����S�iSX����ӌ��6ջi�e$���;1�}�J�־��O�d3b�/��uv������16כ�e�Eߡռ����2�ѿ3��^���w���l��;S��@�a:��ȵN���Lh}�ޅ���w��e
�tӧ:��Ue=��4����q�6�.�~f�~y-Glf�O#�If4�Ph�PT��3�&�t�c�E女�v�׵�)�j$l���W�ZW�6f��r��ů1��+�t�|��B�q���?�x>��� �j�� 7�ՖթN��S��r��w���Ѩ�P��
?9��{�!�<���(�K�I|��tj�qc�Z�:?h��BhK�=�A8�պ�rP�VY�1<�;��K����0���Aod��o��m�	.e���kp�I�
<���?r�M ��3��!W�i痬�ބ���a�8)�/g���rW��׆I�T���� ���(���wp���W���
�q���+�����n��gt�#�E��,L�Y<a�h���Fzc�d��7���N|�Q�&�����M�`�zϴl�Ice9Y*^d�7{���IN�y�F�ܤn�I���IFa��.B4q/<��P��g���|���jӎ�����2�5o�-^����_2D�հM�b�HGad���)|�2�7��үd|��-=�
a+�ţҺ�*-��I��cǉl���+����Z2d�7z=�ؠ��'
�P;_˯�Cf$-_�'8T}:���nHg�K�:���(��v�w�{����(��E*O::
�73K7����a��L�~�<�����zi���]�En�d�N�����U-�"�V�
��orm�����q�,���櫓��)?�Xhpp�Z�ﱅJ��+�Z�.�#Yǩ����d��lj�t������Ǡ@�x�j�-�q�^���ѡ2����͠ Yد���c�o�Ҳ��S$�������������N��M�A��g［����}�k�j�.�k��m�3���o�PL� �荾��;�H�'�o�Z��t��e
�@&�4:�%�=�h�vR��s�_|�g TF��8��������'�3�xk�.���`����}��?F��>"#*x5�����C[�a��o0z��!y���o]��w���=�@v8*�
���dJ��-�
GދV��9)�Z���k-	^Ge>LA���%X�rq�����,�ٹ�^W!���VX|�2�gx���cMG���wi��P'!���^�\��#d�����k8�u�j�w�Uß܊��ϧ"u3�)~.��(h
����nQ��T���p�6T|�K�d����7#�%�ٶ�P�^��|�0zFgd�sY#ѪຐQ�k�x\�Y��\��l�8gZ;X�JO�}�Y�M������:����rk�k�Q�t2���w�C�n�.���p�e������j�O/e+с_����Ưc�+tU*�ٱM��8iL*C���n��	����d�"Uy$��P�a�1��p��I�t�:�g���g�a<#��d
�Ic��&}�i���zsj긗� � �����$���Y�f*v�=@ѕ;��[U�tl	(8�.T��P+8��ʮ�V���w�i�o
}b�%�h�a���%o�H�9Ѥ�9=�J��8�6�U^��3˷�8�^�Z�5s'�F����4��l��=��I}P�`ם����g��g�~)�|��y~�?ɨ���ġ�#�^�µ�����M�r��'|�[K�fV����iTp{K�8��GQ��
OA4����Zq��|fY<̃/e'm��<7��%h���v:��f���ӎ�vᙎ�Uƪ���l������n��P U�Ԭ;]��5���I��,�����8e��p���0.�g�I[��/'<�%��1�\b��-zI�+d�^��p��/~�->�{��IOW�%�7q�������O��}�N8?�*-⷟p~n��_�e7Һ} .=�Q|�tc���-�4���O������x�y�#×U�p�u���S?����X@��+�?���)��r�.>�2�A�&yVy�L�P9q1���?��Ҷ��%}��W�k[�l��$q��z��8U@. ����)��ѹ�&�;��7v3��Fnx?��ItR��'ߎ'k�n��(?��+n�O��5~��f	�Z>t׮tې�ϥS�m�ԙ�7�ON���~��v�y1��H��ҝ/�ޟ�U���$P&>������f���К1��M�YkU�^��j�I��`p��p��N�Q��\��L��+�3~���r�3�e�r�+�9����[�D��q)���B��0�C7��'G�4|��棜�]7�.HF�pv��Ŭ����(�'3�IU�2:�1rN��g�+�h���;�b](<Α�܅l޽|���@Q���K�NF:��.��K�ԙͣ��C��ٍ��T��Jy:�TL�L�#����%��H��4�fT*��3���wO����о|�389�q{��wͼ_��M�)�4h/�QH�t��ecr���,����pM\a��N��GG`��1ΧB��C���KA̟�܍¿�,�d�;�s9Ǩ�x3cB�Iws/��t(t��W�Ȍ��_��t���S�6��5q�c{�:w�Ӱ���QN;"+X�B��N�Y�'fF�|���o�{��o���A����|�sSz�q*�gs*���_}#�9]�HS��`p�WeB�	�y��?�����D�d���,I`�����Fk�K��8y��p��ޅU[�����Ʀ_<�e��V|y���]Tz����4���O�P����Ƈrc>`�x�9�5t*�c�'�8����W���_�<�3�����A*�;��y�����=��D�|N��?�/�7�N!�ڢe���Z��]��B_�g�z���o3��Y��-.<p�;2���4k�?��oy�ۃ��1i����7/�l�Ǳ#��\@��i޻,��Q Ф��5ټ�:�,��m3swRَz`������g)��d٥˽�+�t���>��p��[�![GU){��A�C����i�HF�����'-�&>�u:�3��7Z/mO�����쇛C�t>��kp�����I���i.�K��[��<t>,{��F���ɋ~�H{��Vڇ�A���7�>�p94bp�W�p�����g0'���s�O��GU6���KU&('��T�d�"˟@i;���j���L�J�&e˔G9F�4zrA�Nf���$x���I��5���=�v�2ᤧ#��N���!>:%[�}{:m�N��o��^��	L*?���c�ӧ��*3��ڠ�fl�{����!��qN��8��M�d6�@�=)�2I�{s;)���K����bf�n��������_�R�_�\���R�˟������%�3�(��+����l����z��%�q��m�2�Y&
����(*���9���k�^~���H�Ɣ�-��7���[Z`��ڰ��q
_0q�h`�~k{m�~M�:ow�c@6�pF���1�
�i]t�o>�>~��Ap���_f�N���#�ª
�e���-G�oݥ�����<\Z�ċ��I�
_�ߑcO�������0Jk�t��~�B"�-{�&˴`���x��u]�X�GWA�4�df��E�|􅏓t�NOSHE���v�����o����]4���N0/��F�N&n�f���A���g�n8y��*�.lp{�_���>4����`�O�����s��E�3�&�H�95��%odшO��ϒ.��N���V�	g����,ؼ��?z���|~���A�?V?�[8��3�������8`�z�gh��w���������)z�d�"M���ܕ�+�xF��PM��G�y�7<W~OX��/��t����ֻ� VG]pp��֋�e:�	c޹�S��ɄS��$z����oF��M���w��iw�]���&���A#�f)sӰ�C;4�h����r��wF�?<A^��oa��5K;����-4&�F��m�>5��y�r/:��ğ�+=���En</���R~s���Nx8����߁h�W�
}#�sy���l$K��X~}C6|�̓&��)�-I�|6������XʻcU�kz�WM�N+�*�[��_8�a��K)��Si�߉�ߤ�Y��ؔ��}p�Am�(S�.���&�q3h�����K���$3��Su�ϸ⏎�Hi�w2�Gȉ���Af��[ym/����^�v.�-�~����C-�����R���6Z_��:n�F<:�,Û�c�������(�����<a��|�^��d����շj��5���~�g+O�Kh˦���L��a:WZq?)��m�7-�,sj{�딡��<��f��U�sx�+������O��с|��,-�����}�J:�d0��E�ǝ;��8���Ge��?e��J�S�H$3���Q��c$m�N��Zaj�{ĕ-B�1�����c��1������_8�K�,��iN��HO5TB㑛z3"�I�4{c�)P]���t�F�����ڰ�Q���I�s9�*��I�f�M����хLօ����4n�^�,�K{��c�5"�_�8���9��
�\n3]`Gg⡥h�=B�ݬ�ژ.�ɒ
��utW�.狯�+ѷt��[�1b���o�킬G�ws�T���1��S���3���w~CWظ�T��l�'���ݸ�;�=|��c�m
S3#�L�7��.�xW�,Y��Zk����~���-���y��^9#����lW�\�~3w,�P�ӎLp�n����ؙ8�x��e˻x��⿖kxǡ�ѥ�������>���k��0�=O��V�%�8z��T�
Te��'� Ǟ�a�N�ա�d<����Ŭ����O���|c0±�m��tg�x�z:��O�0��=��j[E��QL<i�wl���:�7a��K\�}�������,�,�́�&�F�E{pp�B��Zs���-�4E'e�,3�]��٦������r֏_N�.e��l~�FΥA�{x^|��tI_�:������S�N�����ί;7���?g69����k�B���~9p�ד��o	*Xs�R4S~�[h�`tύ�������\V_/��)���cb�<Y���F���^�m��}�#1O2�-|fؔ�N�>_�N������B?F`��<��/.�����	-zF�k9�rX���kd��/��K�1�#��S�W3��_~�S;x[�	/��W2Z�+��\�+-�V�)s�\>���Ӱ��e��B��J������x9J��y����W�Ly�<�M:���tV,�����0`���SF޻���؇:c�g��np����{��b��=�<r�]�,��x�k�%jC�x���{�T~�T���K|V�\um��L�2а�E9oV�/z�)��C�xz����^�t��R4��[zE>�\����3��ͩ#�RL{����Zf�ҹ�y�>�̟�Eb)יB�J%����ى�f�OOׯ1R�����{a���a���+6;��k�dV �Rqj\�`���1x'��1�3��+��SQd��̄w���к��F��E��vo�~
��TD-ts���H� fYT��
�я�<� �3F�x��Y���0��n��w�O��r�\e�E��4��54:f��e��]*7�:=�T�K�r���Է��aog�H�
�>�A�e�����4�N��=��%�Ǎ^��O����uvp�U���
���d3SxHGO�I:�t<��o�!Q���Gg�.z񌍭aj	�*��N&N:D�J;��8[�s�^ݴ|�^��DNO���loh�{4���M�ž&\4������'Ӗ��[�{��~�v'~!Zp	>�{�8��sptE�q��q��I��F���������W����%���\�^~��ȱ����K/����l: 3r*�8z`k�HZ������?rN�_��/�'�m�o�pN�uZ(��Q���ִ����6�5~�'nm���	;�`�2���,�:H�����,I�c	O��W��M7%i���wdJ��������-\+XaE�_���Ѧ�	/��F�%��$ރeIߥ�C�E3���G|GT7�N��{Ə2�m��:��t�[��zc<y�<�\k���"n���ދ�Y�<��ݪ��Up�Ѳ��4�-����>����̷��_�/^��މ���ʞ�A0S��pY�#�f᠋jd'�I����Kw�w��rxx�k�U̳�o����A?;E�#�p<V��eM/h��s���2����Lܽe&���6�2�-yG�e���:�ܙN�%V&�gɱux��q}�2��R�0��I;�!q=�1v0� ���O�����;�7Z���ԭ�>W-�Zl����O�?9��H�I�8E&夲P�5��)�a��������d-@J_�ot#=��4u���������7�/��Zt�+N���ɩ��3F���O?���g�p���(�y(����K�Ԑ��hO�VTY��v�=�(l��3|��G��w����Pܻ���.��#�#eOvr�i�D~���_<<��T��ۯG�W�;']+,Ω�]'����l ��RJ�32�r���ȁ��ꂻ�m�K:��� �3W
*x+z�'7�����Cm4R��[?|�x���[p��>��^:\h,	j2p��꘩p8�j�xUX4��7�L�m����d�t��-�YnV'#���v����~7�B-�A�3���i�.řL�څ�wxW7�}/bnq��0g������p{�ZWBS�M6�����%��m/i(�t*�:5�@s���p�>����-��d�҄�wʄ��S�*'F?]�u�^żZ��Q������Y�����3tG?+o֓�� G��L*�>�T# BE�Tt�׶�וaJ��p?�B~�f2@��.y�\���V���s.���U��l':0�Z~]��hk�j37{�ł\�l�Mz�y�'|hL:�7:}	���ȣ��!�9�*bpn�˷}w��1�~�Z_ܨ?ډ_�����)tR~�R#��(:\�,�:�����=<�.����3���?x������07��Z60�n�>�5���0q��z��xa��oxa�2D�F�}O�����tв��^�8��q:1�z����u���a��Zv��;15��Pe6~ԗfC�Y�4s���*Y��o����_��O�w�%|���z��ĥON39�nn�W����q��I6X[ѡ%��&OO�~����ϽR�0�W�w��%F�!��t�Sl��W��e}�,>��Fn��ڏJ8����R�����Q��̊^��c��}2J?u�K_i7u��R,�A���;���h	�g=)�
���5a����?<pc��<�J�4��(�𔘱-��Ĝu�.-��~B#��(B�QH�AҲN'�q��x��b��r�dɜ�����hsoi+���{���zV<���J�ws��{ｗ����${�",��\�rR7�@}�ɯ~��:S_!����xg��k�l�0<�P�=�2���6d��`mBsz�`=[�,
Z��18��@<�AA��M�֍��!h�&��ǇYvE
=�m��n�7�˝�B�¤?;�i2R�hXO& �Q"�n�v�>ó�ȉ��@X��]d-��?�Sb~�TFY`�qF�B�MSapx�O�s�;a)���m�Gg��Z{k��>�NWbs��Дه��$V3���VUߕy����^���^xa�����u������0�=�9e��=���w��Pm���IN�`S�M<:��k��dn���9���	C�h����7�������r��r�w������1փ��� {��F� ���:���.����-ݸ��/���|6J��LNG����ͼ����wh��o�^`�� �&��̷F<����
�]�r��D�����1I��/���E��CKηd:^\)c�?~���/7K.�����)U���^�7�G�����[�^a��^�g�S��,7q��4ǩ�n�zW}�����Ω�T����F�2z'�r�4qI���E�����i�K3}n.��S~
�g`�7�%��$��+�����Ы��_05���6��;��w����YYܸZ��������m��o��
�kҝ^Ɖocf��-^6�2*I��������v9|��:��w���L��o�r9z��
�|��\�CSc[�c�L�7�������~������9i�:��ڔ�o��_�b��_<m���i6�X��|�%�p��ǫ�V���s��h`R�"%\œ.trt�(3�N��)�i��ҳu��eP�Fi�xI��ƫr(ԛϱ��Ə)�l�?�����O�8r�G��rk��P�V�~��3��1�n㞈5���d;�wt'���5X�Y�m9�,y��3x_�g�#G�4������6���7��P3q�f���38j���5Z���+�ܝa��߇�>ѕ�<�\�	BY���n|���CT��wGߞq�������k��Y�?��om^z�X��w���(C��e�VS����d���(;!��_"�h+�e'��Fl�
�ƨR؉2Pu�Y�9����g�����S���	�(�ɪCa�N��e�~��Z��Q���~�ɤ���w/B�#��b�n�Lǃ��E\"�	1
$��YgG��s�ی �>���!7�1�7x�S�WC�?���;y&��;�P�p�y��C����IxR��#�BϬB�K>�t��J/�x,�)����K�=|�������'��q�\�WF��d,������Ƈ��=��2'؁8�y�8��Ϩ~�n�hF��#�����>=�X�q�Me�*���3q�6X���r`G�	�͟��j�f�[h�.��o��/q�����w��а���1�Y��<��qd���4h�Dn����C���4K�O��':4 �pnM>���'߈��cT5��x��M�Q�e�K���E�\U�KstRnyY�1�;~#WǕ6�4�Ȧ1I��S8KƖol'�i��Xn~�c�C6�p���=�ZG���	��_~t�����;�K�׿�4�5t4���DGj��msH�JC5�j?�=3'�/�XZgr5�pLP9,Ë�|	U�2���"��BҮ"$�"����)��&,F�3���6�ƥA�vk=���?|��^e^��?>\�3����yw��_���}m��H�ÚAOz���H9M��%z<N:HA��fNy��X�4���\�>������κrhO㓟��ړG�?���'nb����CxF��;+�J��I$�.�w��:�X�)�w2��/��!߻�%����U��/H�ߍ�J���O�B�>ejPoyd+:k������?�vUV��~�A�Ô9�
�٧�mrr�V.I���q����短#����8jx?t�;�O Z�Eo�X���c��7yG�j�=�P�?v�����W_y�䠵��TWY�m�A=:IO\"�x�	vB��[Ѕ{~������}N['|xƱIi��'.��z�_��6kF0�w"�^H9a���:�K�t�����Ђ�Ѫ:,:?xu������*r��㻵|��?DG��md"��q�����nlz2���/=׃5��<��$�H�n��aS� L�TÖ�1�����K����_z��Q�`+�$V�J̣�6$�=Q�m�ԸQڧh��^*!yd��5�!�Hꨰ��ĥC�ʰ���(���2:��=u��ҳ�_�YW8|�6}�x��FLOߍdӓQ�������>x�����Q�Q��Ѻ�����S�cZ��ŉ�Y;{(<����"�هrxԗ.M|=v<�y^�S��W�*�Ъ�����2=��r͈���3�+S׸��)�R��1:��L�EmSx�w`�Zԁ�gp�۲�5Ht(��LK��R,���[q��� k\�~]�/�Y����k�U-2����^��yx�]�c3~��|Ŷ��(�ݐXz����Gx�"n�҆ǩx����(����72��GCz��ySˏ��+���/��&.y�/��-~��+C�I�Օg�rz���añ������0&n��r���P˿�Ͱ�k��C�Ӽ7_��4�k��"���+�x��.������G�֝83qh�g��O�p�m�3�4��穸eg}8	�3��`�=s��g�v�ѱ4�џ�����F�;���g��RNy_�?a~�o}/�P��C&�#�oq�#4~����[�h��a2��|�	��_=�M�΃�)M���k��ؔ��;�r ?�[..�A�J�ؘc���:��c�r��������k7{��@�O��
�C=H��i��E~����i�on��C�/�-��t�!�Sv7G��-�bs����b�M�e�:��/�W){����nf+J������I+KIN���tYR�6Ѻ�nɨv���GY>���q'��-w2�{���<�Ԓp2�P�s.���h�f,�����p�RϢtz��Y(8���0�m���%/�Q\�x9��X<������(��s���L�3q|/�.�l8!S�{�V]��>�� �؋95I�B^��f�t��-�J�Zz
��Г��K�SoѼ%M��Qfi/Z���8I�`@޽�>��L��֗����r/����k��S�nE.�{�1�M�m{7s����t�����B�([FK�o��/�m�~7K�^}�9Һ���\"��6��ϬAs��6�r�/U��ҡAYna�;�}�a�S�$���޵._9�\��7�>�:�G9}��#��B� OƂ�o*1���^<#.¹��ln}r;��dyK�\O�:�,k�gc��x'g��v�"ٰ3ph��C��8S�����ʵ3P�Н!<��:9i��z���$wc�}�_( �9�+�봐T8
;�L��ȴF7����(�_4�S�_���/?�\f�F֣�ߴ�q�j<ړ6zEC<��e��3M�0T(r����Yt!�� \��bY�_�4Fc�r�͓�����L8Thٌ�"���<��vC�_�-#y�M6����5���1685����N�ǻ�i�6���M���]�y�cal���������%��-��M}��gi���w�&�Ξk�٘u��=�[pv��.��$�b���I�p[|�3|N��w��)}M�@�x��u<���~�?��&�o��[N>Z�.�V�=g��iFy����<��o�#��o䶴��*����#�5����k��w�k^��z���>� �m!68�c��k)�ѓ!���c䠱S�F�l�H7��t��<N���yZ��g{������SN�qSv�<FK����({�����:�}�7�!��4#��>�=�m@=���o�?&p�~}gH����*��o� ���wi�ぃg�Ky;��X������k$xɟk�����04避N�og�i�[�E�)����{d���Ъ�Գ�����.	6a?E��N���E��6eؽ�.#�7�=�Bd�$Ƒ��o���>U����vo�D�~�"�I��P�Kt���!����c:4�15���t�?I�9~a:Ƨ���������=�PD����Qt��'w�Ck����p�qtQ|�N��_�>�����2��AW��0�~k��=иv��ͽ,�V�>����崕�ou��8x�3gT�$�=�iA�]��/�ww33�*��Ic�p'���,�9w��p5K�rH̓48��1��q��+۠������,�z;:H���R������_6)k��1���jOܺ��9���r���t�Wzz��`i	��F��@<Q��
;I�.T��UZ�<��:�.t=̩�
o�^�xws�΍jX���/�s����\x�դV�Oy�L]���yt?{~���~�Nt�q�-?����uI�΋��;�3iP�^>Y:���e����m�}xss�^.0L $@ۿL���2C��~�P���@���>'��C���۾r9���w(!�PKCuz�F`�1xJ��� #Ui�Ͽ
 �5���9Cr�,w�L��i���b��t�;��ȯǨ|�d��m�ß_��E��;l���޽�s����j��_Ǟ��:�ӧ�����G�����:�K���)YK���gH%�����^4��::'-:%���]��nlƨ���ő߸�4F�B�y9~��]�H�O�t�j7k��_���F&`� �K:'  @ IDAT/k���tF�_��/�K���=��C+m�-���lq�l\O�o���~=Ï���~l�
Å'�x���t�C:��o�HS��0Es��{ �U`s��6Χ\�Ŗ}���q�I�,��Or�C��ul<y�du�Ңc�lU�Zf8Ƭ�$�F�b��ю��� �8�u^�Q�ī���w�x��w��>0����gFR�0�u���c�Mo�ת�A_d�������;0��L��B�?'m������Z��qEg����xt5x6ܖ^�8�8iLwe�K��dK�h�Lz�5����Q�#|p��ε���|�k����1�A@9���H�C��$鴅o�O5g��)�|�+�S8N������G�qd�����@t
�����>4�wx6���5^:}��[�/��7<xǃ���e��l�X�"�|�f�9��VK��`yıt��$D���Y�Cn�����N����b�oY��R>8���qaX��{�w�<���9��6r"��;�[�wFS\��~����2�{�w�%g�݌��=�����8\Vi'��=]�����p^�/�Q��05K1 ~��=�o����.�T/e�\��v�ͬ^�0���~�7�������'-����$C4��:n�h=�Y6~���r�h������}��DS�P��s>��n]����u��:����)�KqU�U_%]�
����Ӂ����N:s7j��ًg��\}��P��]x���yk��;�Ա��n�
s��Y�!��O���ŏw�ӽl򿛳Ӕ�\.3��O�M������7�d\2���A6�2 #��2���M���0)�Mp�2�Q�2�$2|�#�]7dF�	�
�U���9
��a#���,����G���C���)�@�
�
�hß�_֠2z���t?�,��K"[���x�����ǒIB�=K�"�e�)��+�ʑw3�_mX�O����>)]q�����F�C<~���=}���m�XC{*k8�r��<Rˢ�UT��P*K|j��u�[�Щoz s*'p�������RQMx�j�u��-8�g��T-��M^��q�k�F7[<	�����ԋ�ھ��G�S����҃-|���4{���W2.r�R�ӌ�<�'|+[��Zթ�$l=��CQ��4�x�ȃg:T��h��FN���C/\�,���;�|ۇ�#��Zgwk������j�;�~�r_����]x�x�w��䦛����u���Y�/�N��w���_�!�Q���?�myCт$pdu�2�R:�����x-�p7���V��G�6~��Q&|�-�k�YZ�H$1��������؝߱W��_��O���#�/��Z��4�P�r�\��:�f�{���.;���nt�wxk�c^f�^m��a�c�58*nt^0O��5<T���c���IS��?a���7'��/n��3x�s����]��Zڛ}}��o�8���y��=�L~�|���,��o���{!�eSѳ��u�I���=̲R|�u�C����)7��V-^4��y�/_�Ϛ���$���������s���%�W|8V:����[�\��ܼՍ�9)HY�]d��m��D#�t��ϝ�5}�L���N�'��8zH[<8��ڒ��"��L��R93ُe�/���ac���ͱ�C�ő�G1|u t�C�W�t��kݴ~�C:³�p�?��3��	� ��ٝ[׫�0�ᤛ�^�>���f(�]Oc������#m0��wA)��'��5���Y6�\�&����˹��Jx�����,I��w2j�B:��bǿ��כ��u2����c��gzmY篰?7<�ݻ:�>�e쯿�Zt�e�g巇2�h)EA/�(Yc1��Yq�F�Q,f'G��$���,ݣ�6?wcl�N!W߉'�í����n�����6���ɨ���o2�����x����l����4og���׆�g(�?��4��u���𓡛�6`�`p��g:A��{Y9�k��*���io;G��v¹�1K�����
G�(�Bw�w�K`�y؉[̈4����IO~�����t��oxY���6��/��o��~J��R:��0qZa~V��p?^��?xZ�a�4�3��w�7�{6ݕͧg�:��
vp*	���'��ĭ�E�$j�_�V��B<�9�j4YjT�yF�����Zz;�}����]8Z[^� �-��E��z�+2
��+�Y;�	#]������Y�1η�9vt�����30�O�#�8��7�.M�����̤Y�[��������;3#��d����<�5\�X�M2N�b�Р�?��g:�>�1~��E;�=�~�/kaB>y��g���5�ѣ���%-�����,[yڭÇ��3�FSX�=��Fd���%���(����q�gu��z����}���^��78���y�!��ͻ:��3:�\���r��I#3��<�Н��k�k������F��$o6���Ə��^5|��/n}Zf0�K��t����=2��Y�,�Z�|g��վ�On��ܼu���K˸����d��:>a��q��}�\�[���g`�es�"%����܆�\������26��+������
���gp,e��?�Ȑ�ә�h�%�w�,���Z��)'�R�S�$)���Y�V^
��.��$M��}�[���y&�!�hN�s��68�M���}i�^����7ެ����7�<��+ ,�{~�ɋ~��ڠ76�.<T��z����=w1�wB/K�r���W�6���������������^�RB/��Cuc���ʙ����\�ג'ya6�����������b�w����Phj@La0B�g���.��8:3���N���iu��P)-�֦i��:�h1�Zc6H+��H�o�oï(C�U�w1�y]8���gf"W�Υ�402j���v���8��[����T�c��l4�mѤP�pPz���#����7�Ə���ptoӪu��)j\����-���.ҨFf�j/�
����
z��;��ex����݅��p\*-����q�� ńǲ�unǌ����ih�m����	w��0�t�4z*A"�� Xt��5�FM�D���SA:�F~Ժۙ������s*>xX��J��/��Ca�{^�E{��m�5����f�H%ʉ�5��=F9��y4ڢC��4gx���ܣ��^ʀ�w�Tz�΋�d3|i@�\ūf����~KG�7
q�I���õVxC�~��٢�*�/mT�fZ?��p��7qɣ# ��o��h�����ͯ.�L��C1eؑe�ķ�a�'7~F��6g�7|)���^Bqr���I�gt��Ggh�i�V�/�K2������|�g�s��\�V�Nx�W��e�\�٥�%�,4�Y;�W��O��3n�������c2	���G|��g�4x��p|��i�e�N�|�:d#���5��n������� ڝ,Rv��\�=-���|�G�����45���=z�_�!?8y�\�k)���Z�ЮeAxH����8{�FB����n
N�gt��i]O����ׁ�C-�'�2���z�����gʤ���3%��#�<k�?���|�{���;23�(�ΰP�E�4ǌ�pN����lʒ�I�x��[~Vu��~N:͝X�2�.�)�mrjfVc�	��ؠ�!$�m�''�W�a�E�����_�\�����T�9"� ~m���4�f�-���^��˟�)Ep�:1+�Ӂx�eW��f��ܼ����w!+i.=�y��/���������MF���or������[�B�gc�������v��<I\
�N����)l�8��	!L_1t4=�b�ޟ6�I$�����Q��'GӒA���
e��/z]~l~n�{R����:#]����W'�O`�s����{-wH|*p[/1PF�5���|����Y8V� �����m��Fc��3�D�∿w���������x�f�����UF�?s��J��8O��8���[Y_i�m�k�*n��h~�����z��S�-X�l6�><+�ubj>�eC�E8Z
8�w��c[���J�e	�X�<�����g�'�o�h��j{�?���w�̓�K��k��6��F���vyK'��j"�ĵ�~rhF��;�0�fՆ��Ȗ���T:~��}׬V1����3|z���w� 
D��YK��Lp�4j�i�����p����`�U�"��m^Z��[�ၮ����Q�I[��?��8��>���A�5������lp}�͐ë�:k�� nhϻo��`�?w�^��SQW�լOy,���x���٣6���[}��y��I�)3�:o�)Wk"vV��n�ݵ(g�/,K�}�;F���J���J���D.e���_&�ۻ���X����J~[a	��\��w�`���N��=�������vO�ʬ����&[~#�k����y���}x�j���ذw|����04T�ޛ��a���?4�_��aG~�i��6�ծy�NV.���������N����(4��6�@Iy�CRa?�ԍP��Ko��~||eKS�v�n/ϔV�Z�o�^��}�0��Ya�ɇ5S�o��W=I޺t��<�a�r~3�$�(�C���b���^��
^w��'���kYկs���-Gƫ�b��)�fC�&��ܹ��9��,w��Y�w�����Ɨ6��~��;���>'Q��@6�z���G��LL�2���ܝ�$����b����ejf7yĽ�[f������##=�G~�a�|7��������V:�W�����߶�����EKd����?�(~t�Y3���TAH��	=��:���5fx�M���rpM|�2s�}�����$8�2��{����R�]�ch�/؂�wd8M�����,Y�~���wm���@/v�#W���G�m�M>�X$6J����F���Rq�b2V�b6.�
�[�?��$�Z%o Fn �U�L��4�X����aF�<ъF?�,��
�Q���^�o&��
�p��*�A��Xg]�'�+ނ_��U�w�;~��9�"���?q����B�,2M6Ua��y9� t��.!J�=�������[�W0h{�'��.�;�p���'�B:F���18��	Vûdc�,�낄7�lY���'qk�?��F���=X�#����?��򫣃�Ī����-��c�x���O6i�!�~'L�8�8ynޅ�f�f�<Fb9���?�%}蚿��D9�#^����-�b'�G�9�O�Nq����{���|�w�
?��I�ږF����3�fOz�o�ލ}��H��h�>g����\9bb����9v��8dk�eKwp���������T�Wl���\Lvח�o�{.�Y�UU��Rn	�r�ѷz�!> M�p�1��o�	��E`�_>h�8�1X���J&���vX���[���Am��/޵�G/B�(wZ�/���,x�Tѣ;uO���iw\э/C��I
12��l`����Dp�K���=.i�22�����܌K��7�8�+�ϫ�d��6��x���'Ҿ#+���%w.��#�&�|�vU��e���I�eA� ��ռ�T>���c��E/�۾lu#eu����Ʊ�뜗@��;��Ç|t%� �n�G/�7x����@�~��AD/o���ȯ^�+L��Ae�E��]#�6=�om]}�Y2�Tw5�ԅ*`�����g�ҿ�^�٫Ư�)&&,*yqB���/��5]�Y�=ܑ>��y���m����W��C{F�>\߹�:t���ͯ�ȯ���N�Q=#^�z����ԙӦ���;���:ۯ�ҳ��o��=yf8��N=з��̆���E1��N��[��.'���0�͞��4�gy�/'9�oO\�pA�6u���R���S��|[u��Ĕ���=�'uB�y3۞���wR�gޕN�T8�\����'`H�JC���y�F���kL,r2Z�R�(>Є�8%���:�t�,��P�ޮ��ˊ��Z���Љ$!�B2������������������T)>&ve��Վ��e*��6P&��<�'�;��d4��H���q􏐢#���h�G9(� ?<�ٵ�l�k���J���Doץ:5� ��&@��O����v�C~��@����_U#L��_�	�z�:�YP�R���C��T�<o�r�z����k٠�.�q�'��LB��9#F'����0a�,p����8�S�o��'3[fX8D�e��v`���.:��	���x9)�k6񖧞nn�q��c�a��|b��-����yQ��q$��o�0&z���,���K�'��×��i$�PSj�R+^��}�R<�>�	�r���B�<�Y����j�[���^MD�Ds�0>�'ϸ};I����E��74��O�k����&ڠ��<��[�K�Ծ�t�e���#z�&)���@s'���p��?��-���/�1!�Jl�<9�Yߨ�C�Ph9�O��|�s���U�mj��Ė:h��uJ���	=e��j?�/2��|���-S��q�>���#m\!:��M��XP;�_m��n���o<���)ig���i�#[*lG��Ȳ~�Ƀ�uVY�t[�\�h4�(�`�aj��Yr���� ŭ&U"��m�pb��?wdZ:�.�U��S!w���m�������ǌ�zw�xl���>���A�"O ����,4Xt���-x��ę����@As����a+�/ׅ�;�%ƻ�@j�u�uU�Ö,
��]x;s�^Y{Ho;:�~H��B�׳Ʋ⅝������~�]�i��l;����7�m��\�����>������	��<crTm���[ú�f�NX`�@�Z?8�ֶ$��l�[���_|3����qU��9�r�5�w�o������7/�z���c�LoC���o��N�(�����H��/�6p�bn@{����c���V��{n+��`�~5!�Nc��q�08����-����\��vA�]I�1+F��3�b�����`I5�V�j���ߊ�.��h�0�o��P-�5�S�/ �J�m}|�n���*��&R;����9�ՉY_6�¶��$���t|Om�W�J�n����ןq>��:����d�+��c/]�ۏ�X�H!��]�7??�iLg�K�a�p/J��/��§l��e�
�uҾ_�}� .~����;�Fw�M ��ke�A�}����:*6r��f`�/�Z�J;�|<�K�b�f�dh�	8�L�p��҈��Q��^i�{��J��H��N�`<tͼ�����4p�Au�z%+����A�#zDv�K��/��i~�-yIS�Gg츧��w�������n�;�����@�0����L�<�WWg����>��<{�]����hS;�=�\zϻ��@]�7(�67?�њ'z& \T�ɉ��[�����ԇ�Mm"w���"�M�N�ʊ�<&��&-L<��V��[��j�����M��d��� ��i��w!�ϗ�Ky�,~���1��\c��I�\�/;b3��ۦX�J]�Cג�=��[�5�j\D?�}!�h��cx3�q]Z��+��|&j��1��O}S8\�d1�����|�1�A.S��]���kM$�>����h�G0�&&�6�7L�"[)KQ��	��#�S���%mё'o��Y8����4��o�a���z���7vCd��у<��mm�����m��uѐs�����=�@�Tb1͇�J�GJ|Qy�!\vRN�Kx��M"HyDq�7����		��W��%��[`�7l�/��m_��z���H�z>�ꆼqx&��[b!�$�r���jc��N�dK��s="�t���<�e,���t�}7�.���i���}�zX��|�����}��1!����?-�E�6<��P9!>w穐љ�_��kQzP������<-m/m��yC�/R_�W[�� ��=-�\`������JVocrC �_&�7��z�7���3p��C�/��[�D��Ę�8�%y��-}џ��X+]�I9W�\��U+�諭��=�_t��፭�^�E94i��q���0����	m�х`8� ����O��Y�5=����&������K���UW�~t��@h�G�+�t����
�ޗAC>� ��K�r.# �Qၮ����{�Km�� �I��*�?lo� #��QF�z�=^�Sp������ɱ��?r��M��~�a/�Q�0т��X'����#��'��啮���x�n�[t��,�"��U|B�x?��I��d�L�LEJ��3t��OxN�c{�ק{��ӆ��x?>iw�q�f�����qBo��S�ph�Z����/<�N�&f�c@��4{�KL�m ݗ�N9��J?&�o
�m6h�+##|�Ga�c�T=�>����I�Ӌ]&���tSr�AYa��������x�lŖ�;�l�HAc^�<:�2c�q��������[���S�i/�#_��
�r�tb>���ɺ�g��S:M7���ցg��#���%:�#L��l�`m�0	����񢌶<~y6A萣�	��K�>0�9bl�/q�;ədC��$\�x1y\XՄ4t��~|9h��	�N���4ܱ�y�V�Gb� y\>c����@�� ���=x�G�����.&�]���K�!�7�/�ʇf����\�Hsd���S����t�(7�&8�=y:/P�x1	�F����-�����kh�o�n�!q�F6��%m@��3�w���O>�wn��c�� .io}�C6�/0.Vs��81�zh��U�!�����:�.��p�܌�e�N��z�G��]���#K����� w����2���|���.pЍ:x�0��C�.�#��v�`�_��s���k����	�)z�����ƶ�����H���O����t�l	�	��{�#��T�Y��]��	Z�S��Ï�M�n��]�3bxQ���S|��Ϡ�U�*5��crgW#W8bf~j^.�;�����#`tH�D���'f�8�F�<v34}0OxQQ~�\
�&�e��t�_�J^�|^�\���e��r�r�tߠA���r�k�~��U�uM�~�8���o?��AO{�ksC�,�r�M��T�+��7�hZ�>/Q�VU�cxROJU<^7XY��*t����cLo����G�m��4���Zދ��v�������o����l����_��8c�(�%�:<B�Y� jo�x�������������n���n�W2Ŀ�YP�+i�Y$T@������t��ޞ������S���+ ��%��R)����C��w��Cʺ��1��<[3�h`�g�����p�^�h��J�;� ���L؍�}��|��`�k8ɉ���.�Sѩ��4m����;���M\�F�����> -q����ç��?��Ի�}���<{��w�ۆ���7Ui�eAA�|_�]oo��,L^31*=��߹�����fѾŜ[�X���[V�x� oL��¢9�_L�)!.z����U��^�n��b�H��Oh�i Y�	^��H����>^��]}���^�JzGs5���l�&��i�ЄGt&^đO�K۞ӑGwh�t�Z������RW��E9?$`&��z~� ���{�8��8�zܴC�Ñst�8r���y\l���"}�E9���&��g�]���Nשq��ޱ�3/�)�@��-AV�R}"��<3�B�4��Zxz:�j�x�O���>8�k�Ƃb� �PzR�~8�����q^&�8�
��8�%�֗c
|�x�<Y�ϲ�8�Q��F��N2�#��[;p���z�UC��Ɇ���q�ˆʏ2�ʕl��-�"7�����z�,b{A�0N������K�f0B�~b��9�Ϗ��
�hp�'��r�)c��=��N�j�uGy`��&t�x�:��M�	��L�q�2�48��GEi��Ѧ-��9<-Um\������ER��91ȽN�����E�_{^��I/���e"�#r��Gz&Z�_��,1��I��4���jh#�C�xӥ���	�7<���O*u��E ��D.�O~���5�Iàtu�k��ۆ���R���;��;�V���Snx'���<�F��Vz)X����!�'i�<B��dX�wO|���=m��&��y��S-qd�M&y��i���0� ~�Qm���Q1z�"��^/�򵕺�_���*y�bR�$�=Ҝkя	��q�W��s�cC����&�`đ~=�Ď:��"���P՟葟z�<�:�~��<Gd4w���uy��	�#M�<!>�"ƈ����v4?�|��6B���!uI �/�CH~Ҕӏ��>e����K���g�ܩ����'?�o�y��I]DGd˷\�����o����I��s�����@���?��-p�{�/B�]�>�Jp����Ne�Uj[ϟ�����I��b[��ll����!
������%��Ä:��|�ы9�b�ړ.$��1�x�[]�ofy���z�GF�9ʒ��h�=��H�3���D0r�O/8
���xt|0H�Z�֪�.s���[�w�Aw�����:�N���d@cY�4U�+4m��~F��@��������=�I���y��
݀h����Ą��[(�xh(�j��D���JÅ��+VS���"$��i\�<��ľ蜸����)E-5
.A�VV���)�89�C���z�Q����ĳ�i;�o��|p#���9�)�ş�'�l����������o6i1FaJ|�L6uiܦ򁹎�Z�>D���XmDiY5�:ŏn�BSe�6N�^+_W���a}�i�	օ՝%Pz��&�/���>_������q���/	s�{>��yh⡉�pЭ ڵ��	e�/j��c���u}�/�GOb�@���dO��|לp,&�Q�]��{��F��^2J
����|c_�L| G�-���O`���w?Y)���wF4�pyc�Q=��%�]XQ|=��$�7�c|�6��v�#/��o�?����s�w�K˫mA�I��"?��_�G�2��9�?ᔽ�/��!E-�/_2�-��@K^�uA�!���gC���c�7��ŏ�	/xd�S�zsa14������?�5хg���N8�\�}0	Ϥr�OdE614Y���9O�/4�(C&��˳R;z�����{'�K;%���+W��[h�/�gŵ5	Y�F����M�Ё�E��@��;5�꧔�N�}��yMs�Є_�H��[�x�ݣ?��l�cz��Ŧ���F�r�BK�$��O=N/����Gf��y�A!�g�����y�-�P_����䓽�zI	��W҄�)�S9���O�����my9�V!A8�����R���'�� N��aIS?*�J%&���x��<0/��«ZT�b;�&���*u]�S�w-���ld0�'��ѵ��|�)���L�P���|�����,!��R�:b����c����AV�u�n����o�e���Oh���.{���P���E6��J��x��:R�I�&m�U����� 9Ĭ�����&#?q��=����.�_҉AA������s�G��������v-?�?��<d��=��yl^����/�)�=�n��A���D�	bʍ�xGF��GEn���ÆǢ�vO`�E��f]yq�7�~x�&��1�Þ���7�X�Ɗ>e{�O���ͻ�L+��kL�.�!�0?�� ��/����N�'�2F; 8�8h�x��V��3�%O���p�K�\|��
������#���s��3y|���I}HY�ЀX��k���ѷ�/����l�=�3�!?�_�|x-�ra���}�r��2� ރ==��1�'v�'����/���8�{��M�9nW�G��������8|�N��j2Y���M�^���҆�{�HB�	l��k`����&�*�",��/�O�q��A�	�,@����}�����'�	����+�ȃ&�xrׄx��B�g��s豋����`{��������r'�4:p���;LL��C��9Ѐ�����K�O9$�X�$�v�r�3�љ<|S�y�l�|it�߽Œk� �T/�Q]��1�u�2�`<��O�@v�}8�|I=6<jn��W!�   ��M��TN F��	�IC�S�<	�1`�ɡ�n���"�<���^�z5e<C���u�i<i�����E�Ĕ3a�ib\ޱ���Q�
lA?p��W  #�n�O���&�L�`�c=HN`��(�kQQ�	L��s��Wq�Y�&�����)��I�V� ^h����nt���)�c�Xeh�)f�ǀ�eS%�!l��mI{X�����Q�ޓ���cң���pqO�a�Gz�@�
�LL̻������ ���[K%5	m��R|k4��ӝR��H[��F��k�c�>���jFS1�ԅ��\5);G5�������&�6���*M9�_�7 <zח�G@�n�>g���˵�v��`SF���`:��-A��(���ӌhz�=��z�F�1�-�X�V���p�b�3�o��0�ixB.�[�(+J�3��#��UA(�>m�V%��5۬����5���ݣ�,>K�IN��h�-_�}�F�#����wp���.���o�P?�<�O�����9���z4U�����}��I]�"x�;R�_L��C/xƇ�o�c�|�X
�,�Q��Й�Xu�蜸���4|��[��[��|��p?��O_ϗ��ϴwI.b�Lm��z���h�)�	���K|�8<������/�pL�C��/w�Ʌ����ٝ}��_��P-|�x�7���pg����,��ztb��g>BG�dS>�<x���2If��Ŗ��^�����;��V=���/�{�Э�MC�ݍ�ՠE�����v�X�;6�y>`mcM��C~6�x�&�$�����<�5N���:�՟n;��ėv8׮�����ڶ��z�hM��ɿh�o.��Г<��
��A��@�
�x��n|O|y��n�W�"b�D=p��	�`3�Ya#1/Xx�R�����yyU:��!?i��6�-O��Ox�bt����eh��ǹ�q81�aൌ��"����_������Ž*��Kų?�`�Z�!\�}�ᤡ#�?i�i�� �*;��#`�~�~��~�^3�|���o>j�.�Bρ��؄�s����	^���,1��L�>&M9GO<!W�9�y᫘I��t��	��m�2`����^�a��^��!O�~O}`�g�֘C�Xpw�>?�n_o���e�H�7����o`��
n�.n���G{k���Ge�����|��-9��7*]D�w�O\F��ԙ
�I!�����O@�O��m����M0L�z���Ӣpj��I�B=��,Gi����oB�IG7�ԡ�2] ���0.Zsi}�w�|��|�6b��8a�Uߓ�^������2h���P΁�Ĝ�z^��c;����تc�`"e	��y��x����^�3�Oƃ໏5~[�Ϟ/<	=� �����#	4������fph���N�Iz7���qe=<{\ҁE^�S|�X�qF��2<���*����yv|�#2G"%�?ʒ�<:�6e�e�<��zh��0����礡#$-ǥ��4�:� k���=ix����#�ւ`Y��O^�z�)]�[�+S��꺾qh�x���������}��g�Ο?�t�w�ygx��wݗ�{�9�a���W������z0�={fx�g�U�Þ�gR��'�,�״b��z��ɽ���`�~��������_��_-�o\�����}���韆��������_4�:���~Q�k��6�;wΓr&�ׯ_�x��O?��^�{�oD�z�����W�'N�:ߪ���?���{��o�S߄z����?�����k�7��xM1[�V�-�#GK�g�cǎ�z����B���xF
~o]��P�i�i��QZa�J[ޏ�6�[���j)Ɏ�^mk_��
�VSh��9����jw�o^��ւm�㤴��'�=uzX=��[I����W�.�]��0��{��]tO'�a�,����ک�9�pSo0Ъ[8j5v��TF����`+���;�
��[�y4��"ֵ��bˎn�2-�� [m�Ӫ�Vx���:�`UɟlWc��C;T��{�@���V�zrJ2��;{7�^bt��,�ϞE�u��А�����~!<�6���LP'be��$�ܼ���ٛ<ӶQ�CjK�6~c���0>�@���L��"B���*��''H�Z��_�vդ倻.�/��	�ސ
��Z����;Ʋ�&L�����S�%\U
W���̬��:�
����犩Z�����bJ�E�ֽ�˕_�u96� �j8�dwᩆ�o�
?���cㅼ�6�
X� ?�?���-��B���eq/�i�j7��(��T4� ��fI�:?X���]B��W�	�K~ʉ3o3���[w�A�&ɵ��E��¢�?�!�\�
>��+8MW�?�����a;Ү��^�����T\��C5\e��8��M���uE��[���,���)�������~�Ki�m�eF�h ��G$���Β�"�M1֍c�j�WJ�ÎGF�0��x>����Ԕ?�0�1��\�p^r)�H������D�[����%*4�(���DטdK�y�,';*c����Ho���-������C.���$���|�ف��\q����6W�h���/��G�ÔQ��,�6���/�%_�ӯ�UN(���0�[��s�k�0�΅4��(W�A.�i�N����z���eFG+;��ߑ񂶳�*�th�CdƯ������s�S��vB���}�Kt'._ɷ:gTz����s���������}�y�T�������[Bʝ�r��?�����%���'_�RڟvƫUG��꒽򜚙���}	��&/:���A.!��;'��{y��uNg"{�����ן��p�����SO���_\�^x�O��Ϥ���C�����? ����3�/z��_�����	����勗��O=9|���M}0�s�^}�_���|�w�==�~`s��|V4_ἂ��������_��_�;ځ��ŧ�ѻ��7<q�����x�W���S��x����ցq��������[׳g�j���p������_��cs����o�GW�q�x�����"����ҒbO��O�\=|y��?O�>1����^�ܐO�ᗿ�]�ض�z����V�5��j��:�9\8f��̥�g�Ν9�݁a]cݒ����P�?����׮��U�Ǐ��WB�>�zK�/�\���z;w'�#�)�Σ��Q���iy��퇶�6��u�`p�A���k6�$l�k`���ؖ�|X���Uʩ��)}��������2���DR�/�ޒ���VH_W>��eՔ��2qc�ML�r�(8�ô�S�<0@�Gp���d��e���)� #�	8����FV��d	���
=pb�Ǵ�O`)�ea#�����#G��.�)'M�w4}�7�{\���&򔥜���;��_(.�#�<��y+O��^-���[Q�G�LSL?����KF_�t�CtOY���	���#yʦ/IO~o<���+��4uu�;6g���l�)�	�rO0AZ��M���C�C�J��Z�t��>N:xH7����Č�� 0@Ͽ��5|e�|n,�~��O�����|1�g�}�z� ��M�	\r�&�t�=��	��C��?t�x\^œ>Ф,����uU���:Г��8 ����Ѕ�8�L�U�<�|ÃA �Ұ��o�?�!��<�Q��@�����-�;���d�g�g��Wmbx$M�#p�)xBp������9����?]}�).������{#k�/8�����c?:?�=�B��|����c��m��M�_b  @ IDAT��"�(9��gސ@�����ᕮ���h���2���C84^T���ޒ���K�n��:L�3q%���/����Lp!������U�˗/\��n ���b�@��7��#��}��{��;y�w�x�M��w��hxU��Kw$����9����W[������e����t��O~���W5p��+��U���K/�4�ɟ��m���k���p��3ß��?ӂ�o��o��?�xx��-}��֝���gL��G���_{!�W^���-r�`;���������>��9���oex����rڶ\����?>��}Ѽ*>�=}}��D����Z�pх/�S�{������g./������KÙ�'�zX|Ew,�B�o�{���چh�6�H�Cñ��O�~9<������}�mP�ۚ�j!"�iԥ֧v��T�o���p�%��5?hof��wue����������O����g���W��0�Iv�M̂bUWhͪ�������_o������X�n��54c��v&xӁs��fz�����8h�����'�N�_I��ٟ���:,�8��G@e�C/i��u�bK�ph�\�a+�ూ�v��~��lO<��|�W0����&Y����@���Ox�Rxth���I�x��G^pJ�i��d]Wy{�Gh�`�1�-'��ǖ� ��/��-*j-��Յ�i�|�ȇ*|���`�S���?��c����7�����o��K����N�l1��#l���"T�ҲKi1р7Xu��9~Ѕ���X'�����ej!�l�C��8}�<��Ӣu��	�ۡƑ��|�7�b��t0�O�qPz���e���,i��j4�8������	�Bk�r��(��k1H�A��X6>���E �V2S��S�ҹ��H��t�C��_=^���6iU�+�3�{Z���H�UtaG�٣>*�CU!���J�/���nv��b�2���t�3BlL<��'�<���C���dDo�H	��O�]�*hҫ�(�|�r~3Q�	�\��?���FVOc�ν�t��=�e+|�At ��ad_;��"?8��;:��غ�������}|��� ���0�tp�:����"���̅8¿��?�<ґ��S�VP�֕k?���~��!Mto���zw���yqp��i�������pT[q��9���w��ӏ�O�ĉc���L�?���Ë����:�w_�C��w7�]�6p���^Є���ʻ��_y{عso��ؔM���=/N���3�ٸ6ܺ][�����p���W���p��������䅳ަu����W�zs����Aoy�!�;ë�}�w-^Q��?�1\����'_n�8�I��.����ݶN����bN�:1���׽u�l;r���_}���a=�mb�tw��'���o�Z�\�"���/������.����L;ز���<��eZT]~��p�̉a]��-�X�m�9�7==��$�+���6��G������kñ�G4��]������.#��]]����^\�������&:DM�=ig����2Q�`Mȏ�6��˧u��8wl8��-"6t{nc����1��a����!=���wb8�=eO�?����?�3���zX�;�es	yl���#���^�SwV���{ ��,(�lESi9t�!��O�����6.bx��,�T�#�G����P?�`�9Vg�P���1B�	>YQ��	}:�o����=�s����>��%M��Y���"��UO�=,iʠM. n���
y��'G�p���J�cq���q�Y�F�^�}��*]�<<B3YV����	:h�sp�4��BnŤ��Ȫ.�˗EC�6���l�3_����h������ǎQ��w�w�M�-ۋS+3}jj�D6�Q'���|���A���hH�.g}�/|�=��v�m�����)�s^��A���?t�3i�>��1�D�,((��n;����l)!�G�Y�	��%�8�E��f��'��;�:4����L�����
�2nST�BxW<���pxC��x��62����,�CV߆CKy��a��d$���$�=:�y�ώ(�����Ga~�o�Gn�����#��)#��r��ܹ��	�����C>��%�t�ZbB�>�Ì����:�hwʣ8����܂���������]5gK�
M���p�'��|p��G�L/Յb�j��y���C9��e@�>0炖�؁W2�"�����Kl���n��1�&�j~YTܽ{{`1rJ[�,��5�F?�s���'�F��.?��ǎ[~;u��`ɶ$�&�<u�wWxF��;x&�O?1��G�[�^֝��t���ߴ�l����W����}'O�n�����1�᰾�9\�/>�g�O^�|Iwq^��,�n���۷���c\����]G����O����^|n8�E6^?�b�����c�ޭ�iԟf�[K���#��!I�ҡv����no�sm�y[ݗ��V��y; �vc����jpNu8�}�lM�����N?����>=�?ǳZ9���cJҭ�#r��b�ߏ�O�2�p�p�Yת�Y�`�z%��g/�}���w�t�i�CC�-Q�j@˃&T�4N%wȣ/N ��ah�t�
u�S'#��	S88��B��=�䳘�3���8>�)��|Y���ϑI��N�&���I ����7���<qp�}�9d�п'�r&q��Dξ1�ξ��G&��3O�sC��
6�pR�	�ʪ�[|��rœ��]���ڂ�/�?�
��������8��<龼O'1e=pë��ҋ��}w1A���U����Ap�粰/nN*�ډ�lf�!�
;Xg�LF�Ș�;�=�jҷ�����q�8��=���C]�唥ϒ�/��>�/�ewG�eB��>��t�h:Ʉ�Ĝpz�����]����/C,�!Gډo�BXe�.���ɠ�ߧv�K����[�A���ɖ�Љz��-X?��Y��Uҧ#�o��/y��u��w98Ҁ��<~��4��~|Fľ�^�?�C�-؎ۚ�#/�u�LH�M�C�'x�}��RAu �ŠSo�1#B7�{�/sj
 �q��a�)�C�#/�߾o��	]�	��S��18�'oÕ/eI�yA�=^�7��O��]������G<�G��E�>�j���c��lpC,Gt�� N���`	�A����踟��{���y�[o��m;x{[����H��o3ag+��Ç��Nj"�;\����ռR/*rZSF���ੋOk�x���6u�8[}��v%,.Ё9ϧT���D�����?��?���������z�8�	��Q���?����7�gU�<��/��?,�n��~�������x��ޫ��n\�P;pn�!�-�����0��;<������aw�-�v�0c����b���G�W^}yx��g}7��u�\��s�[�ӓ>���J����S�st���p��ԅy=�̶�������W�,�q;�����o��[��3GNc������N2</�����@��W_Փ��y���9u�	��$9��v'n�C=��Q5�`-�%x��Zn�Ɩ'�ܩP�H&�R�Rx&���&�4$��1ѰXP�gO9��<�y���#v<� 7q�l�B�������ӥ��W8����%f����-R�Zy��� �j�߼�
OB:;��8�D&1<�G�w���"�'9��x�����	m����\b`9B��\L>����fۏ��'m��ğ|��|%��d[pC?"<"�������ǆ�ʀ�}�u!��ܥm���~���%��~���!�Y@�}߽Q{a����\�`��o�(A�(!\d��@�-a�iħ줬�§����iW�R
'u�x^�*-x��ǁO��+r��GYB�@BC�<-	��� +��'>5�I��	U1�|k��E����)�g�����=N��qt��y���*��|�!�lR��k��?���C�����NĒ��L54�E��g�h��Y��m���X����o��kc�vx�oۤ)c��S�6G?`�M���n�[y�$�.����
���<������|���%��a{�'�����q��Ĕ�W��hpD\�;?�_o������Eq7��%�Àz��q��z���q4-yʘ�0�eN��S_V��Tz W���܇�s���g�/�����e�/}^�2gc.u���aUw�h��Ǟ8��*��je����m�zA��O�y���sO<1<s�Y?S{���*r8�g�u��q=D����� �7������Ow������A4�����������m���=�����״��ysw ��C�7�7�P���t�w���W�������<�>\��m9�><q欟�`"��{���L�A��_]��w��h�'�/�]鎾#���y���o����K�h���p���}��wp~����<����'W�3Z|?yzX�B���^�V�-�y�b��.���(���nꃋ�,s�e}�C�ˡ����J�	����.�!��9��i_߸-�o���z�Es��ke�����E����*oY�mi8��Q=U~HO�k���^�z�������|R��U��;���nO�j�\��G��/'O���}���	t�a�I�e��1j�����dF��#��t`L�y�a[ogʂ�}�|	����(�h4t8��_W�xRƊ7�޻�b �ī�k���N��r�9tV�5-*�N!rH�S6x(Ml�tp)��s���Iy��L��
_`�'��=�1h��1�ʉ�'P�ɳ�N>��긎�� n����nz��+��y;�*���S�b=���\�4B�jOo��D�io���i���~����9n�X�NŢ 텖�� � 	�m�pR�^���zC�?&Q�X>P =ϊ��$�l{��K8W��窷H�C�x�u>��+�,��N��M|��Ƿ|̱6�?P��JkШ:�4�B(7���h+�����Җ��G=C�Ў:��ԶTl ���2�E���TLz������n󅨍�b �;r�66�I�|���zp���ӛ�Bo?���ͯ���O�z9�R��$L��7c7o�b{0ڐL#������;���2�[��sl	���6VT��̠���~�&b�z�,�BO�h�,�pR�B��>��lg�τ�7�5C2�@K`�+�o�E�{��Wv���ip�K\��~x%^�k#}�'���j�
����d��w�hux⢪_`9L#�~�F|8�g�;�/��E��,(�^�3�`���vy<pԋ
��c^�w���0_���1���A?�,JxF��J�>i�����-��z��)m:�oܼ}W_���>>�:�y���=�L��+��י��������s�->�<4�B�ҥ�^t��O��ݻ�ܶ=Оy^���?ԛ�^��[�wGi�f�����&�z�&��6�&����MM������>��ß�9��ß���=|������s-8������+7~���������&�g�,�/@�9�����k=���_�V$�r{W~�+�����W/��~u�����+�l��
X2��=� ������ᖾL����w[���^��cs'Ϟ�C����O��uxNo���z����=�Aϝ;��/R��O'�6�c�/P(�\y��[z���..뙊;���{Ú�������n_|~Sϲ|鷰���?�0o�~�]�bʭ1�5@�na=u��+���p��I�*/h/�a���d^��o�v�� �A�[' ��R4b:�<��չvO� �t��)>�CQ��*F��#��t�8^eSudʑML'� ��NL��������=��M�����-��ˇ��o�_Bx/k!G���-~�û��Ӗ�*B�)��6t���`�e�����|�]�CI����+|�A���B�� �u��̱�p���(�ѣ����>��8��q��\��<�$�A�,��`�<���G���j��1z�`JY�'Z-	M����4,7����T|'_�P��;d��Z&r�v����.{Zt��|hL��=��MY�Os{��%��a�?��a��`�9/C�Ȧ��}�/�S���aI�|Co�ޗ�	�z��BO����V�t	ܯV����ӃO`B.e��nC��FxU}N�=]p̤��Qli~����h�,i�TXP�\�a�!Z�`�]k�:Q]��Wk ��a>�?}>�l�\l�͉SV
�Oй&m5�e�H]Ok:���gl�	q��j_Fj?�O\8��7S��z�R�đ)�q��I܄F:�)'���]�x"(={��kr��Y w�5�� �,G+v�ÒN�}��S�Ҵ��Q��ȼ8�$&���c"�E�zU?s4��Ib��YXTp1�yNB舱��b����"]�Wt#�"o�<�~���ug��=�?�������[>oy��ϥ�/(x�2nܺ�I8c{��w�G�4c7������Um�'l<r����έۺ�pe�������G�hP���)_:�y�����x�Ï?2.���]�Y�.�䛯���Gw/�j�4>~���|���ulM����}_~v�w*.\xj��	>ob����B��P\����3���g������������z(���������6���G2�̺�Ʃ�޻��;�
������������wu��Z��vն�l�Fb�DmM���C�:k�=m�Z�\�+O'��^�t������õu�������o�U-\9Tʞ�,>�m�%5�3G��מ>9��ӗ���1���*���n�=�^�X�r5R�ԏMՁ8qzl�*J�񠾨H�?��֊wE���W��0|��'��Mݢ{xO��!n�=�bj�q���&���6���:,�����%�*Zֶ�ϯ��ݎ��Mu�e9��,r�:"�b���Nt���diE�tO�R�4�͍��;z=L4i�S�����x�P[������*�iuX>I/�W�+j����+{t��z舫��&	����'�~��.����R5��[��J> �Ua郑
0���+]�`�v5�֦љ�zm>���'�i���vF��C���T���B�D���2���XV[L �7�t�"_���%C�t��z$���+������>��NW�֑J�Bo�e�����E��/�bBm9Q�+���ϸ�T[�DE?#K�Y��\�H[���A�׀�t�Ǻ���`�_�L�&yꐷ蠠�)��<k�d���ܣO�?�1m���C��%.P�FÐ]�Ǥ>#-+%�:~� �[V%]xm�i]��t��p����L���W�_LA���-H#�.�2���m���Y��T�ˆ=��؀#޾r,���� 58����8ا��&b�+�a|Dʊ����@�yőU0�-m.�7ϒ`>�#��0&���X���J��
����f��b��l�x�G�歴mu���·��Q�u�ζ.��+wGi�2��^�����]U7 Fz�}�@&��k��������zb�]w�2y���H�W���:m~}+,u|�`�����i�5)e��[���l>a۹�q��� �,��-����Gt��_�s�ץ�HP�<c�ht%�mK��0^�1_Zpˆjӫ\�K.�xk:�W�|��	[�r�@ȅ$�M~�O��J��hŃ%%tmxj��O��L��g�Ú�*�#��XO������x����o��-u��B[k�XLr<)�\ z��Ú�>�;��2͗�e�d� =���-ջ�~eD�/���&_}���"��\N'0ݙ�- ���U��1�Q�n�=�����tH�i���`�[m����EF� �v�K]5ߖ�z���#�~��59��0��g�ϯ^~7���l-���;çZ�`o|�=�5�1�<�X���T?��t�R��l�bW>�X�ƨg,8�C{���a������m�9��[w�_�ï�+o_�ݙ#úvذ[C��&������B�"��߿eݢ������v�`��o�j!���A? 3YQ�<��y�75�5���n�)�	�#m�>�����C���;�����J�oc[�U�;��Z>�g)�j�2�9yH)=���Eh��EoZ6��g����> \��\�ズO�tNɠ^P%�9}B�HNˉ51Њ���`x��(�좃5A#FL ��qh08���U�������MO�)á���͇!cU?78��[��_�����s�k�����'ÿ콯]� D>t��Mf� T��z�
�2%�L���3�%^=~| /�7�L:e���I�@�;1�I`��#������=Ab�P�,x�1�����B�Г�,��p��'���3}��|S��	!��E�|bp������OF�s��YV����hrL��3r{}���o���e���s�=���34��OΤ�)�m��� ^/�t�k��7?����G��wES6 ��G�N���n� �bt
]m���~�1��`j�`0�3�p����:�{��]�C1ۮ��@�ڷ��b2ȳ='p�!�`KAt Nڌ��N�=i�80�h:�4�e�%N9�#cX���X��~j3���8�|��1r����/8��	��Y:=��/���⨋�6Zx�N�7�3����I��+�n	��&��?0�����*>~N ����"�\�>�v�����3x$Pf���՗%��$�t*̔%�lɛ��"�䷾;��=M҅��wr.W_���<�h�Ox��B�ű�Kk���D��e����>�~�Q��������h��`.E��.�_��C<���6�~�@�&�a���w�i�,7�z�R7���$�s���� �b�|/���=�m��'�� k?H&��M�H[�2&���>���]���#�A˖^d�����Pʐ����A�ޗ�H{���4wF8���v[�A�q�k�٩�[;7�zٛ#�$ ��~�歅��7r�����=}��z��x�1�٫�QϺ����9��ۮ���;)�t�����)�����ߟ㣡��,��QscEÐuH�}}�>�ws�uU�\:�ձ�"��.�m����y�l�+�x˱8�+!ć�xz@g���{�K�
ƕ9�B��=���>]���:��d]�Ʈj�At{G��!����胾�s�K�,�aE�F�+�M���ɱn�w��p�;M�vvJwb�$[mo�{=�s��x���?��S�8e�����2��l�c��ӧ��T�?�'7䅷80����)�v��ى�X�km�L�CF�O٘�7c|�i�@�	݂@R$dR��>?х��_�Sh����7�}���~Dz��p��$���.��3ȇw�7}����-���g��p�͠~B�#0�'[&�n���L䏍���o��mI�/�q�۸cl�\(#�;��+��1�x������'bл�#���<i�1�ڔ����S��`��>+�(pw1�m-�7��6x�S�R�x��>�,��%Z��~DG�s ����h�R���|�P2������^�	�����yb ���d��pN!��:�G|o�~x=���C�����v�'$&|`��e�$,8��q՜+���i[�݈��Ȋ�ģ��?��F��}O]x�k]�*��'2�ǂ�~
I����҉W䀏\��i�*��s�/�}������'�g��"�r���k��op�3�R*�x��� ��8{xY�b�mx����f��}�7 }r��2/(4��q՞�5 xo�U��YW��o��y�s|+��2�����d��=:3I'F?�U
V��bi�H�P�M�q�e�ǪQ��)�s�R�~V?粗�+�3u��:bQ /l�v�`���/<{���ȸ��8�}��=�B���i��s���&�[��Ȱͼ��t���zS�	�M=F@�r��AՖ�A�m�Aχ�������� 
�`�跴[�g;����ֵѿ�#����y���U-2ure˃N�jh��j��G���u9A��-[�����������n��I����@Q�	?iCǹ�°�x����xV�^�cC��u[��g�����;'��`U��{��Cu��Ձ�芐�4nd��U=V�s$ +G�K�����fc�|�-rh�i��Żh�W�J�����%M�/rn�w�����Ѱ�>�cY;vv�<�n9��]cl@��-u�8�9�5�z�@kT`�ǹ���m�p�1�#���k�Vj���9_
��-�AV�NZxQ���3���|��'��8���u�6F���CC��wE�=.8}���l&ܦ���G_*î�AxM��C�H�CC_$f�g?,'�\�`�7NFlu��/d�Cq�i?S���Bח%-�,˸�N���u��4r�x�/�b���N:�Qy�_�W`��Sn ���<0|0��ꃲ�I�6�#��1r����b��CN���dL�����i��I����ׁq���:Mb�H:2�	ё4<L̓����t�.�9���4џ������ke������U�3կq%j�7yxrq��q����� wގ#���7a�P���BS�3kށ�B�"���~�����@��{ߕM���$�/�ybW�i�,20N�o�9R�?�e�-�	��0O��,N8�����V��==ߪk�5���&�����41�XPxQ�q9�҄�a~�I�\g�S�ޢ�>t�Cy0�1y�}R�����M�$�xm>�).��5�����������K9��Hc�a]0>\,Lώ��C:z{+�h�}(����ji��;�����lY���(oߵ�/�����WTt}���I=��I	d�m6�ѣ�9*�z�wK�rq=gP�갇�^W����jiK۝5H7�դ��a(�@
��D�S��
�6����miU������+zG+B*w�ɡe��VŏEϲt��7�����mlj�����Fb�k���]!�ї��A��Hű%�4�sU���ǫ@�J�<yxi(�^ʍ�~�Ѕ}����n^!�&'|#\�lm�*����K��qq�a���*ٝ�y�D�(�nA���W��d�K�E�>�9�������<3£��p�]؄�V^��&��tʬ#�Y`R��zL~#˲[����l���:���W�D��.�11ph��z8e�	}ق}�/������f�������_g�71�5I����
/�-�M����˞~����[����[W�𚬱�Iǒ��g?}Y|1�]��\r�x-Z�����o�m���ɘ�_���S���W�ղe���E.��!0q�W��_ПXlQl���n�ۤ8����_�Yt�&��J>�����Vw����jB��Ռi�K98���1r��~�|�?)�kt�B9>���M���?z'.���Ԧᛲ�{��~e��>��\�hZ=R�?�y��p^*;�*��q#]o��c�dZ�d˼�~i`�	��m� ����@~ҁC�1��Z`��I{y$P���L��E0��Ox����9�g����[���ߐ&�|�<5�Ҥ��&σn�m��Ӡ���
������<
t�O��<|���	<�U^�s�kر�~�;h���<�n��'1��Bg���|���0�{>�����$x�3��JOt7�d�,�Ǣ�>hw�k"\x�'p7�׉���A���<8уtBpl��G�vVʘSFq!��1�)��*�|�]�������?��	�~n(#Mʿm�Y�*C��CT���X�ۙ�����i��rk88�{���[��G9q�P"�c�,�-T�����Ç����T㦳��:�3���@L�)�S�VI��ڹ=l<�w&t��/���=��ӓ������⧓R�8�4@Nա���*0��4V�lI��ã��,x�=
[�����P�3�4�&7e�Md���81[8(ωt|�Bg
��:dE���|G��$�(=���3�+�ӄ��[�z��/���w������>��8�Zq+LYp�{X҉��|�����Q�����'��'��2����)�#�H�8�=�(o���|��B/�|�I��1� S����)!y�^�{c��;ãƃ�f�BؼY�ڂO���z��?��[�������}��&�8ų��Y����g���uM��O>a��׭�R|S��C'�Q`�'qڣ��O��<4���Ȼ��
,��^���8���I ���_S����~	~��!��]B���7�"��	O#�~R�B��/#'px���)�����i�Υ�>�)<`�a��w�%�oB�K�����兆��������^����}�ۚ i�8H�G.qp��.�a8>�v��,ˀ@�t���]��v�6<��4���~	,`|�A����#�x]tt���aa����C�����)}��	���>�~yk��ךC�,�z#��0�%�?Dy�2��$p�#����CK��GW��NO�}��@��<.$g!�OV�B����6'��N�?�ccx���<�Sƕ��)�I���9<ȇ���#�l�
�>r�V,��!f��&q��\P<���Q� t��O8�1��0��<Pw�T�ܡ���U�����c����a�� J�u�3������,4���L�-@�3X�����9�9*�%F�+�N9���(OU�U�� nԺR�/� �ѽ]�Fk{�ΰ��BZy��(נy_oH�}�ְ~����A�L�q2JN@4�y� �o�'6CC��Tz�!�����P�!��)O�6�z�>����,�5�,(ƫ�ܢzl�Z��9��8���-�ߙ~.���5��O��W�K�I�~!�I������#�}h�ƌ\���ׇ�μ��g��]�X�_�ZsSN^i�Gt���w���~�	��}�����#;z�~���f�ͻM@�x�D/y�1�S�ӑ&�L�q�Vԗ)�����6#,U �h¢N�pt�O�\�l��eC�7�(&���+N�et5�~�4�w���ǒ��U�L��-u�[�Ϙ1nӢ�\V�_�@����=�D���	^���ʢw��X���~���7?�3/9ѓL|��G��7������!f��x�+��:GEF���y�����~h��e��>���r�����[��g���4	���	1z���&n��wM�C<Gɡ�Om��4"�2��c��cK�0�����(ph�+}(<��=�<px���ӷ�0�I�E�p��� J��H�q8��f䉎��/z1��;�3'Jyp�'�n�Z2c;t�����sÏ��p��q=H�Ű��eͅ�w�͇�{�Gi��kHy&� ��]��]>�6�_P����C'Bʈc{o�C9�c#4���X0y�۸�:���y�=/���?s��`�L�r,�\`�<B~[���p�
N[E�I��'��$��`8x�`�@��21ꕒ�ͮM?t�s�ڨ\�_���Xw�tB�EgvJ�X*1�&%WM�;V��f'Jg;6�*S��w~��-�KL5`�F
%�Yn����1ހ������w�2w�U����NE[=!3���9(�
��mCoiʛ&0(t8��KH8��0n�S�Zo4��Pܡ��Cٳ�׭�ݾ=�ެۖ�Hb����,��*�G��`����<h	،�c��\:1|�c��ª�e���c���Op���<6�������p�c~����1��G�ѳ�Ԝ�tj�FM��c��w8��^>�<�r�9}�_"O�7~��)��M��W�Dg�r�#��K:p�)����'��	S��2i��9�Geс���F;%P,��ml�,h`,b�! S�yM��s�O�?4ʍ2S�8���R?}� ot�����A�4c	o�L-��WT���G��k�a*�kg���%� ��r��Ů�s��pj0�Ƌ�~�m��vy!�<�ĭz`桱�8�j�Y�(0��>��ɸ�SO�$���\��%B���~�����]d�1p�<1.R��3����s���2;}�K��<|S�9,K�!���R�~�C���
���)(r�ꑼ�+��7Yx�	kt�~M6��i�k����/r�zd'�~&H��@nߏ��U��36�[zb~�7��+����8����9ȣbd�r�s�|Б��"�Ą��ۨ�����n��Ї_�'M�O��Dt��4u<pi�9���u7�C�yLx���ŧ�^~�y/(>�ts�D�q��`a*���9�&�:"99�y���y{�Us��m����N� >� <��>)�WN�)������b�~W9�	�91���1���Fj?��p�/��lx��:�O '!���������=�׉���Py.�|�>[M��v��7[ő��|��~����zh��m9Ff�2�����k-�XW;�x���p��������!9c��M݊���(x�nɨ]=��p��
zB���>��Y���G�
��������~>�{/z�����W6Z�/ZM��h�L��������{�^e>�� j�����V*��&��_�_��F����ō/�]��7膧� ����,�vގ*�&��U�*�����P+�K� �
"��J���U��\<(��9Bg|a�<��777�M�5�qG�a;���.�'ߓ��wal�4�aY�:�y���UI�N"��kk�rc�^�o�U:�+��O��byd�hyP����+�ć�p��.��ceς�<t�/��a[|��.�Q%��f��h�G�MZ�It��ѡ��	�~�F� }�=Ӊ`�M���F*DqtL{�`Fibʢ: �r=<m���8|��a���2@#�|�Wݦ�]r�~ヴ�5ɿ{���Ln����CMp�:�|t�L]]�W?�k=�>m���@�9��sp��̣��:�"���5�
�#c����؞x�:�� L*�>���R Z������
!�ؾFG�����N�u[d�Q�?�Q�)�[�]z6�С�����I�[@��6!�\"��m| 84�\���	d�XX;XwUB>0� m���q%r���*/�>l�Ҧs��d���+��%w�YT���{�ۆ��`C��a�N*����c�_�GZ�-��z��pY/�༔>/����Z�3����F{:Y�/�ɏL�yƴ���kY����es�dԷ7�\�n��<K�hȨ����mCu���9��]���ó�����EM���j=���T�YFK�퀤�c_>Q��FuWVV��d_MU=�χ9�G4}��� K��yKN{0�:�\�H"|t���m�AWڇ���?H�����wgO�gz�O�h4��	r@�H#�a)��.t�?�Gx��x$�� ���������zΩ�� ��Q�c�}u�2��s���RWK/7)D�d���!��"�Z��h^H~�3i�q_��=G؛�W��m:��B�=~��Ⱦ�Le�����{x'���9���+�����<�O��Wo�Ʒ�<��Z�s��Px�2ָ��m�+���1��r��,�*ò�O@F������M>����+����++x�shO��Vu��!���O�ғ�t���h\�}�,쾧Hy�z�������MR����,:�K�h��~���}x��/�K�2��_^N��B����������R_};m��o������/_;\��O-$���2G�~z��;����4����c��7r��zg��&��ѣ6��O�g���B[�Q�����?���ʏ^�L�������':��94��?�����9��y*E�=ϩ���p���<I�deo�U����y$d�c;�����|����������L���月�夳�	N��As���y���It�C!-�Ҍ'6�R`S������7���F,�I/��ەE&��-_߫{c�V�ȯ��$�6v1��"��� E��#�')P�aШ�#un���;� �c.'%1����Z�Vh4V(?+#̮���Ƿ�;��=���XJ�R0Vծ��:U�ڛ��ROS8~!���k�L2��9/��/��g��ƚF�E��Y��6�U�5�Fh�E*6#�Yv��U+-�U5V���"V&[�kń�,G��b÷�WG��Iq�}�걆٩���&-E�/��z��}�[\���K�Aj<�L��W:+.��?��:��5�E��F�<m�̎V��>�f��U�C������S0y!Ǣu�N����׆9�od2v��|���J��X$7KUS� �_fE�T�C�P�q�� ��^�������Լaȶ�= T�EI�	��Rk�Agׄ��-GEY�pg��'��͌{��f'&��k!�oV*~�t&���y��U���}�~xБ&Ē�$�����GZ�7W�̇�z��YLS�[��*�$�n_�ol�D�4�&%��t���t��f])O6�nW�p�P��-�4ۄhѷN6����ӳ2�I��/�W���}����ͭ=�w9%��KRew`�}�,<R�#�~�f&r~\�V��d��&�0��®"c�|ٴ�
%tBI�K$�x����]�%�]���!}F�R�,1�#G������������I�4L2I�_R���	�)�� m�:lV�z����y0�,Z�-���[���aI�� ���k۹?��$�����%dB<U�H'�����yq��]~���L[-��A��I������:�v��]������[��@�K�Ap���"ˊtB����+�P���َ�2�b���%�����߳�E����j�Ov�� ��]�����:�:�}�^�J�zS2t��x�eg{�F��~���6���\���T�\�Q{�#�S JH�	��Y��� �N2Hpe��Lbd�J?~��~�s�8���0"�fC��	���l*g;q��������k�#�
,�����}���,v��Nr��U��x|��J#���2d�~c��iɯ����/o1����@��)��c
.�U�;ƿ�#	O��|��o�&��������  �s��)�;1��|�D��8���\�)��]��t&ű/�vUb?ʘ�-d0�?l�Yi�ڿ��9�j6�u���g>Gb�������am������(���b���b�9�*��`���h�\?W��p��T@At�l�Б ���ǽ6#B�fk����At�t���k�ҐEaq���|r�=�9�/�C��ݝ$�[<�v�h���2SB;��m9�L����'b���/s'8����J��)J�,r	����!�l �w.��Grn���^�J�̋�]߹��u��?ܨ����;�E���wF��&�����Hx���P�+�0�ɮ��~�ū���r,$Z�~�6Z�'1��VBg%,�f3��U�D�e:��p���I�|��z��VP#t,H_sc��|���2���*%ĸ���Z2�7#$�8��;�Qt �U8��I59]$�FI�1?%K*Z/Hh��| ��7>�<^��u�J�Z3B(v��U�?�^�Jc�K(,���ح����\�ͫi��D�<#�5Z�U���� �X�|���?d/���.��<��ИX�\LVDC��Bg����a!�"�s�䏊�`��|J�?��-p\�lpk��{�v婀�!a%�B=V {�斿���g���l�F�����,9NϪ�_�:�3����l��S�7J{��gI���Y�ӳ���g����,�)��5�ӊ{f�	�&��MrI�8X�tvo�u��(�(�.��K��u��d����%A_��L�t:����J;�%��	�oi�8"��A�L/����Z�ZЀ��Y�?d�_]´��d���pg:�# {�,LDS��G�>��qs�#.Mj�i X`��m&��iD���PZq4Hw��VԂ�%��O�J��έޤw7��B�XnwG.����I�*�e�ǊӖ#��IW�#K=��؁������j����H��G��D�]>Ϯ#���7)OR0%�ÁL�SaU���i�}����hXeq�WG��H�:��2��/�E`� ���K	���ڳe�h(bM(�?{�������7�%	6�|n�8�1;���d�ےb�'��9&�ûv���Qv��N�.��ƽ��䬙�O����JS�+;��R�[;&�0ǡ�:(��(_��8j=�s�����،O�ޛ,� |�s���/r��֐�'�6���H�������B���n2��D}�7�BGM]��6kTל��Lf{���N�$��M���=�MH������ق*'�����iS����i��u��k�~{G_���L��*li�<��\�n`[�*��8����{���Eؼ9����b���i� C�fg���ke"ڵ)����EHH}HŢ����l��āp�|�<����
���sZ[�q&��c�L2�������zB��j���!k_�s~h�X������v�I������A������n�1I��E%f,�;߱o�޻X�R"n{��Tk��u(S5_˗+�j����o$�^���^�?8�2�XZI�B�i��gw�E��M�A�jȗE}?Z��iBoysG{���7��-�y�O�Z\�.�!���]&t9nx1��ag�� ��#r�Gy��Wp�ks-Va>@���Z�Ѝd�g�U�������j���Ŕ>�9`<x��_��>��<x#�����7��2'/#䒜�8�m#j��ߌ՘��W<�a�I�
��M>��Q��T�����m��nx��R��#��2�cE�UWY�Q�t�yPux�=B�v�q���}x8�F�_jb$�)F�=q�bZ�[��s�,�}t�"�D,ds,����$���%0vw��Qҡ`9�V����@����V�˯= MuFA�]�����y���縻[1��	Dw��K����={���eyl�xX���[�ܐ�����&||��I*�6��ͱ<+#}���%��_��u�G��z�[�@9D{ ���ԑj�M�Y3�LcaM/`ӯ�R��ܮL!^��N'�D��=���u�!۟T��6��~NUi����?yw��L���W.���[�����G��~^G��.-N^e�z�Ǻ��3�8:�IΏ�¥A��b�!V�;Q<E����ؗ���,,��4��<5˗����t�T��#�/l=H��#���������\���v�j�g��]l�h|t�[�2"$�!�|�G<�e%��_��\�b!ؤ�s�<�1�I���Z�A�<�����?�G�gHC`���`O!O.��SduP��4h�^��m:�0 ��R��r�g_���{is��~C#�Г��!`	{�hR3IZ�Ovߎ�o�O��p�O*�H23��WP�!MJ�Y[����P������;L��V�t(`���d�OvY��ȓ�)��R���R�Q�t	 }<�6��}h��f��0�5�ʱ>%��.	��i���(@^���>�dw4�%��#Ŵ̶��y6o��H8>�K�!��6E���`.��V��1`a��N�+���� $���5�hz�uOF�"2�_:$WS2��Qk>�![˲G���~;��-x�����Vk�ߑ��SNje������P �	R��|��x��>rƞ�i1����"�t�j����U:���k�%bӫ�b���|}��G�	'��'�>�jC����K�t�*$i�d�p���EX�����k߲�P7�G��Ýb$d�lt 7�&�x<�yy�Z"���S-,{�0Y��!-.T�� �Q&�����Z����K��F��'��3���94R�`����'�5���mHN�j�l��b�&�@b�q������Ϊ��aMz}U
.���ө'���6\��&=���X*~̤���%T�7W�]X��1�������MuK��<Q���mڔO�8=�LDr9&(4�E�0_�,�����\��������[	�rz|',/�<��[�誸���X�-$��K$��j��KѦ`࣓<�R�FVL7����7B(}��
�s�xcu�Z!��2I�B*{������{&s����%䣂̈́=8y������uμnDn^F�pbffէ@B=�����za�m�f)fK[����`WP3<�����MW���%�;�>6T����Vȸҭ�>`S�d(���R��x����l}�WR�����Zq�H�q�|�{#=/�<`�#����]b��x��M�ޜU��?z)�x;>�o5�2����걧їǢ{ <��e��K"��*NO�����Q���_���'�[eb���C8��s���k�ؾ"#Ӭj�w'�;�*_x��$���$����JJ���.̘�f���ȉ!�;�%������hC�;�h�����˕QmH�{i�9?9b�|w���Z��U;� # �zք����Q���us�$pc�%O���m�Cɕmҹue(�J �~�����=���Ţa*(��J��ȹ4�'J.�xy$�Y-D�$��G���;D]L�zR'�b^�z
��ػ<�\���v�䭚��i��<2;�_"?��	�G�o�m���w ���-����Ib�I8�i���r=�ÿ?I '��U8�&QHShGs͍���������_�N��|��0�x�\h�]�m�PJB��L�^�	#.��q)�����x.��u����IE�i������w�_.,�\+�X�<�l��$�y��nX�ٿ������N����2L��k�^c[�i*Q~��/��V1�N.�J�VNIC�a�&=!YL��8:���g �,,���x�"�����f]���U�}Ob���K���ju_	f���f7|�>z��3�._�x���-���D�����@��~iU!p-χ���Oq=n�2S9�!)&>�%�����p�~�wQmc>9P?y�W�Ϲ,o��3����Y~�O ��R�XJ������f\U��[6*�1�RH�,��������B�WV=��lE6�b�2�z��$��b��:_)ko"#M7FK���g}�@g�^�U�~�n�c�9�퇬�?漌l���R�YW^%��vp�w���5�Q���.�,Aps�i�I�!��#5`��cIYֽ�Wq�IM�6P�>�������KI���]�F���ӊ0K\�۷!5}^�aU���ȗ��p=��jޗ���I��6�dv�^iK=��ͫ���J����=1v%�FWM�3�(h$ĥ��D��'0ֻn�v�oj^�찈���ĉJ`h9�\*�ƿ�Ɠ�L?�r��A*��K>A�l���~�z���|�4nQN?�	?*+���z���ҫzv�H��n6����z��	��0� �z#�2^6m<�Fj�V�72����40�;�E��ø7�!)��ssy�4'�qGK�X��PE�B�p�f9 �C����V�k�%\4�ہ��w���/�}�\ʢ��('�5���|0Y!�Lٖ��2�w2�<Cq�����C��?H�-l�G�2��\�����s����c��Μ&�����N����E�]���K�����t�h�G*���C�Lp�!�IQ�?�[)��ut|���+1�~��*&},���^
��Gi����@d@���|'�(��ab�܀�M���6�Wv��e���;{�)|)�n~�a잺O�QJ��t��'|�J�ǡ�^,�t�Pn�����^u��������̰<A���{TmK|JP ���A��2Yl����gL\!��h=� �h�Psd4�N����V��i�tK$�����styq�ٞW<x��P��XH�:�"Ꙍ�J)��D��v�[�ń}�(�~���Vjf1�����3��k�}�H%DH��&���U�k�B:���e�]����S�ù��ͣ�d|і��[4�1y���>�6�աη�d ���$�XS^Q�P&�6{@S�����Pa�ܮx}��RK�������^�4���N�JYu����B�2��wX Чz��O�s�(�yZ����� Mi���/D��3�q�i{7F��=89�6��:بg�6v��l���`[��<� ��}a��{��6�Ѧㆀ��*�޽�LfS��|)�"�(#�4w��+l��T�V�����C�a~�6�M����Mh1�pe �KǢz���h�Ο�z��^؂e�#�k���R�1N։s��lMk�:��L���H��<1mM(:a�+S� �Q+�6�C����ȥ	��=U��+�	��Z�f��o$��ѻ��xA��}�	(�ͬ"����T�z����*?F�2�8.�!�F�^�|���������m���;���L���[�6f�u%[[՘�,G}�Ț�
g�f'�����<.���*��x�_�JK"�� �s��������hh��%���y���B�w+�<��|Tue��sy��!>�#"=);�%�ȌƔ��|��G�.��z2E�Z�RCmo�]�����t��gx?֕�,9s�.��(��-BC(�� ����%���3zw�Vr�$Wy�"��GdP���:<�.<ML�d������y����VH�<u����PiU��L3_��SfZ��c����٢���c,�,�t�bX��|kEڢ�Vbk�i>_wF�Y�y�5Q�'�=���l�-y/B�iL���=E��������ߛ��'>�A��{p��^�����a[ߍ�]㟿�^z����0�0_J�R��Ig�y�m�c���UT:i�r}?�iڶ���)����6b�>�}k����VM��υ�-�etz?-�a��d�{
Y�o�_�tbq%�����w�Eg��Ń�ñ9I?I��R >~}�i�QFB�H8	���^����-��S�*����3��s���/�EOz����*��oO��<#w�i7[�|P^�f둺➖�2!�l,"�\���p�L Hg�"@�F��]/ѪM�`��,Dl��(��R���*��7Ԣ�sv������O���m�r�mpo�'B&����=2B)�K�O�-���d-r�o>a�o���S]\?�jm��Cw +����U�d��եs"�ê��c����z/<e�C�8w��:Owg�����X^���\
ꏉ�����B2�5�ݔ�ݏ��ڰ�1�,apTI.8�s�������=Ko�k�Wn�����Ē:>eG���4,�5w����f���0uF��P2芒���`헀�Yh�C�=�8���l�vx0�;Z<����YԷdx�w�憴��g�s�}�g2�������-D�C%/�D ��}�}�u�Ie�����ꛅ�E���] �E�<����Hfk��o/
������ӟ�zD\4�6j�r<Q甐�o��e�������^���5����};ʏ������+f���W}���8���
�=w� ��	��脧�/���D�~��JƂc�LEC��YR�.�`9ڄo����L�w��ƤWh]'¦N>T��s��I.6���2��� ԡi���=�Ǭt��� \"�&�'�5���f<�x�Y��@A���/�wO}�-�n^��*���,d1�*���Xײ#h��F1g�Z�K��˦����)�W��ϫiD?�ʼ9��G��|�V��V��Z��r��v���<u9@�m�u
ݗl�g-?���ĬW���́�Y8�2BΣ��K@���ٿ��-S���S�c�M����
e�f�f�X��Z8����^��h��c�K���rc��&���������7Z�c-<âwS~W7��v�q��5�h�Ƹ�~�g����_Nt�H�ܿ��y:.-�v	iU]P�[��`M�ł��3+�x�&徰l��ސx�%�@騫ͪ����Us�(���gx\�o����6���Ytx�G-�7B��dkxrf}��'?�|�#�J�`�pIH@}� y�p�w�@�5׹�ޜ�؍FՅ�d�|l�x��۲�������-��-���ٯg����E�wU���~��q�:=y�b����X2\9�u�Io�1��]��f�:��r9�2_U�z5H2'",@���3\�H�,�gQ�'>!x+�B�Ư���,�����W�)z��"��v
r����z���m��ڔ�PBP99�X���_��R�<��ŧ:�G�3O����,�I�d��!˻�j�˲oע$O	>����i��
C%.� ���1�`��^Z��[u4b����p���)N�U���n!Mj����XQ��B�U�������>�O��-��]��Y	)Z�Z��\ֱ�aT;р7�o沇p���-�m~;�P���$J6k�����M_I
�]�]fdo�'�i�m6��0}(���z��G���}Ac[�qˌi�_��[����F�n�����L���(���nvՆX�-���.�Y��x������\#���w \�1҉|A�����n<����K��:i��D���$���Zx[����2@�\=���҉X��\~SDq~���.�	��HR��*~�9\�lO��V���3�j:Ky���u�+�w���q�Z-a�^� ���c����	4���ņ�5[��Y~���vV}��x!cϚ�O�]��	�E���������p�'�V꼎�~fgY �*�`�g�*��ө���~/�E��#�;��
&Z�HHe+��e���jyH.5.;�$J����$�X��L�;����	�@Ur`�Ci�D�.�zq�}1��>�r����Fn)����ߧ�_����M�K���K�p`SZ6~.�Z7�+1�&���H�W�R�=`�ڨL5㼑H�}9��B�V�V�c�}F�;F�0���e�h��qz��o��s~�ĉ�}��:s&ʗ���y%|�~�����d3���f̱>�
p�1�� �"��e��h�����Y
q��R(�9͐�t�c���]p��V)u4&R���	4d�e��r�%0��3���F��7�e^p�%�{w ���8?.�C���DVg�K���%؉P�3����k�4m��D�E��{ڰ/��������Ӫ�B� ���8X�D��K�� ����7���t�+�nW�R��V�"e���f�Gb�tk�v�ڏ�,���5�wy��!�ƨO�@�x������kqf���O�$L��8����y@r|�|��U�y��<���C��;m06��Bڠ��UW�G��i���*�%��q�P{#ѣ���G��}2�i�k[�a"��9��Y;C]R��u��3�K7��B�?rA��	��\�R�H�\������>�-���:��f6Mb>�i�0��vCUљ��2&���'��7�M���UMc��WRNe�3F'�Vc��Ѓ���B��a�oD!��)=s}��vt]�ʥq�-s~o,�Ϳ�rp��KP`d���].|���8�4�?0.X����l�_t�j��iG�8%�$H�J+J�k�|��ۍ���k��.�Zmu伣7Ѳ/l=>�_*u'� \e�A,��}P�X�%
w���5�;s=#��`��
�]��.g���=��S��G���bC��}�ה�,~+�v���(Q�pe�o��ć=�Tt��������T�h��,�f �6U��XIՄ!�{j\Z���ה=$��8S^�C�l���-@��(��Pi��y�s8��.'���^� ����]`�ؐŖ���+T:��H�zc&x�+�ƴ"�t�=+�����ig�ΕR�.�7�S�o��ǝqI�؈��+����Ћ���>�&Z?��K݆ /�<�t��OTa��Y[ �WH�],ol#��e4Nϥ�1W'qS���˷�M�-�_��!�{1q�4��S�4s[R�3 *�T˲�8E������]:��҆�QȖ%8T���j9��n@)��Ď����6��u���&~7|�!��Wq��O4���X|�+j�<:���[�8̀����E�
��)�13��:6���h�F�v-N�n!�/ѻ�
k�������Tu?X�ԠF�;m�n(\ę���~�N��&��#!Y��_�0��S
�AT��s:���̞��Lƚ0��s� o6l�FS��$]l�����/2E4g�BvOec��i$_HT>)��8b)apn�g�>�pY����nM�`A'��h���$��F����`�T|�ҹr�׷^�	8���v�m���Km�q-�B�P9���hp.�]S��n����z:}���;���Lkس<���M�f)��P��k���K}g9:~[8x9�WKm���E�G���	���:�94)nڴ�N���yJ���^p�<��t���Jh�p�v[P	����ITuUXB�U���ܙH�:��-�Hͻ�l�N�����Sy���UT��[�{S7�p��5uaO�<R�UvV��}3�馲�ۡ':��3���]h��ҕg�I��j�8^M���²���0���ó�`���G5.?4s=tMv��r~u�"��^��t�S=|#ئ�	�w�~�X���l�]ۂ}��l���`&�=�3���]5092�U��~ҍ�M���[�9�<W�e����-��Jv���$�l�?+��Uo�Ԥ&'���ʻ��"|��x�@��DO?�^7l�7Q����ٲ���,�Q᭏�[S��J|��-i��aT��wg������U�"���5�}�]�Ct;�Rj~l�Oi9��@�.��r]���;�k4P�����y@�{�C��2�ܰ{�c���ig��
k�&�����nѨyڼ	�o��Պ�^����-]F��LMtܬr(����V����VVo�c5�ڳcfn��3�����e�� �Fb��9{1���}`:i9���h<��������=�³�r�+�ΦCN*���������˨Ea�����י�$R��BKS-�s�����)���ܽ�uW�{�'s|�Kk0uZ�Q�@�̖�{;� �{�3�a����.)���|q�B�W��Β�f�g��c��ܳ0�C�����%7��j��"��o2+���ۤ7y�<?��3^�͌����	�@��{��:5�x���R��q�^-��Ѡ��O���]-K�(fp�U�ӥ�����.�3r�tÿ�U~���'>ND��<���|���כc9/�!�xB��A(x�5����5c��� ���>����a����0�	��@?��n�v�S�ܷ<�tWt7���v����0��E���O�[~���y�g��+�^�_L����VX����
��ҟ���r3�����ߜ�tRޛ�A/eN��h����y������Ė�$E1��`�Y��~d��Q;q(p���$0��ՙõ����?�w���Ӑ�t���8������z�w��x�6*���̮B7�oÁԻI�1�
�sҡ��L|�?�<�Eqku������r6�F�|ӃX�:��	Nu[�^�-b_>>�m�<rn$�ckE�J�'���=��p쫨$�Y�kc<�`����݌MZhidў�2����d�\���r��������4��q�a��ҭ���3���������jm�Z1�\�,vW8{	[���Я��Y�yUsr�(
��V6G��d��|Lq7�Pί�%ŵ���gkU���yr{w��Jt�[�VP=��S��V_~K�4�E�ߞ��>�ܼ��М�|��]ӭ�z�����H�u�d��f<͕z���b��f��ɬ6þE�l��L��ƛ�F���3u�\6��氛kYB�Ϯ�>���L����U�[��u�|����������,�ɼ���5�RU��A���pÞ��}^2��3~�zn'��T���mmZ6T�ߟ�[A����c
���o��	����M��]R��J�ؼ�j�T�Q3���>�6h��c'�����16-.�:wZ%�U�d2�u�~	�n�r��ߟ�K���6����Zc���Q�k��y�~�c�c�T=8�	y�U��{xP���u������'��X�ܸ�&����	?E�(�Y�1�U��	����)��l�};.���2V��V�5���7���A����0��h�^|a��v!���eg�������	��^��=�U,���ű߳�ړP� ���##pic���t)��z�w�~���G����5<���i�����ª��N����T��]!	�<����ӹ6LMh�'��{�6Mm��Iv3)�sI��1���\�Y��*W���q��zj�z�~��f�����8��Ox��d?���")G�9 ��������m�8hӬ�+ C��
�i��RU�/���+�����Y\�y�mz�B�J���M3�<X�u���Ft�|���o�/-֚���߇ɪ&�sdǃ/	�T��i�m�Z������9˯z�>;�������u%X�p��\K�[���ˌvTo�xW�S�پ���ۊDI�ٷ�sB��+��1�ǪO.[����z�ӝe�t������M!��Q�Q(�&ɢ�̓{�_�$22O^}��?���L=ԁo��+3V6m����klvy�@�����ؗI7��Yc���τ ���~L^q�,��H�+���M4H�SUB�9�І��q��_����@�g��W�UƔ��`,��^��D?�̙��{����O��V����[��Cdԣ(Z,�z���v�ak ��Лq7 �jF�,q�1N/Q�.i�Z�q�=u���-���d֗�sE�'�%�y���S ��h�6o�w��S�N���tS���J8nf[�WU���.w�ay��?3����Nw�坧����V�|�?q�2��e��ӆ�\����s��途:��?��28|�{���`� �/-)2W��y'��Ԫz��� ���Q0���+���iu���4|tZL�H�@���Dpyw�j�<H�bP�����E3��lO
=R?[_���4
o��E�rF��,u��~%;��.6��FZ}t�UU�K��Ե)a2��&�i|ˑ>4�{$_��d5�|����w��ȅ�#JlvV؂��Y�b���i֬e`��#ׂ�ˑ�)*�4���Z����pԘ�3y��s�Xb ��vԻ���0'e����c��c<)�h%0�:�K�iٹ;�v7Zkf�z"��@�!<����2!OS�I�w�$�A��d�_�sl�?�7�27���;�C��kv��5\Ү^y�!�Ց�ཧ����'��{�3���"����>�n��&�A-k�~e�(�~�^����"p�;�N|����������R�Yk�u۳����P�����/�����J�/�%�������0�I?�3��1 ��ck�zn&�����,<P5C�q�^�t�N����R7��2��hNki�`'&Qr]�b��C@Z�H�y.t!��~��;C���ڌ�EaC��F0�K��R^7el%iA}�5~<�8��s��y����8�q�J��ΐ�,�Uy�CS�0�O���m�Xc9�:F3۔�7t'B �c�A�g)j���`�g���
^y�Ԗ���{��d��;�=Xt �>�KN�)S*�b��G��Kۆ�S�#Hr�Ƌ:��/�#�ŵ7�,��E�wbt2��!�B?K�v��~,E0�e��m?9z?�#�8rŸ3�>����z1_�SF�����#K͓�K����t]-�i9������B��fu"�'�Iњɳt66h�>x���"��}A�uJ	����F�#޺a�O��^��Ʌ�݅<���j��H[a9(���.�G�~+�����p��ˋ�5��C�'�Z�x���o������)�c��Ni�v	D��7�raPy�N?�*�p��K��-��!��53�zb�4��C��)��Yew/T���.��Q�U��(>[�:[�@�
tZ^+s���4i�^r@h�8J�LО��w�f���G-*�}<)^E�[#����F*�qlӠ�2:�H�!�ٴq��W6<u�m�V��|�K0k�R~�T�]ajI{��r
��f��`��y��߿�ˮ�י��Z���/iƳg*2�e>�E�G$���IU�־C���3����|{���dd/N����5�,�ƛ�}�7]��ZY����7s�����^�S�55��W�7+��TL�d_{d>ӭ��my�,[��H���=u9a��U��)�g��nORuNn�Y��@s��1=��WA��'���!���"�rh��^Cڤ�%��ف�V�㪯���_p/GU��	���|�D�[� =�λq,�T!~��Ľ��t�s>&�z������s8q�������2C�ɬ��=.m7s�2}�����Inq����>	�U}��2�NU*���V�y�]�j��>��̦,Ӭ�u�1���6;E�fE�����ע��z��N�US�r/�ar� �4��3�`�T�l��+�Rސ�Ցs�QS�h�8����:���۶YP�P�Y��yc:��B[t�y^�.O%�]������4�u�r����������]�0��d�f�b#��eQ�ֱ��;M}s_�4.��|mL�=�&-C�y��妴�u7ð������;��Rg=l��rw���b��*�z�P�u6WC�q����B���n�0UQ�%P�zۊ��Ȥ���#��+������zyx��k��5�� �6IT����M���&08�:��Ϋ jQ&/���R]����l���1a����,C��8��<�O�<��N��,E1��?L����\�d���	lr����r翘�Z��TM�,���n�C�P� əlvh���R9�7�4�^酯=�K�\Y8'/��3��H*�5��q�?P�ַua��Ԥ\N���B�i��p��e��:R�'�b���1����K����.$����V:�D6��~�lj��{{{
B����߇���f,�s��6믢�)���8��f�t y�2��p�h�)��W�����,\ϱq����WH��mU	�0QT�^~F��rQSNfy#�E�}f¬ ߰�	��=��e.�پ�͙��z�R8D����4v]8N0]Ϟ�����?�( �/�hz�~�m�bK�i/Y��^%�q�v�z��o��b7�t����F|�w������.N��G��ȟ���P�m��(�������+L��.$hv4_l��$qb��wU,�<���'7VO����Ao0�/ti��]���.'�h��bl���&�O*�%9v��=8��*���^n���� ��l���.��S'ci�F��ʟ�-��[�#��7��X8n��)Ƿ�W�"���+�>ibCv	��\8�7u�J�NfFq��c��i�έ�_;��(~Q�{��WB�����4��?c�v�������{����hGiopPH�הs|.$�ɔ��6l?a�Hɾ�&oO7g1����֣�I�j����3J��,�������������3�:���p�}r.�+����V
[�p��q�'\�@�S����� ���R��i����3\��Tɂ�*���uO���2���b��J���[�:B�&&Q���XF�918B��9��8����,9�_Z�2���-J|"��r{�	�1!|�cͻpӄ��(�D-y��Qf�;��'��n�]l���f�Cg+þO�{]Dɒ���J��s
x�z+��T��6����k�X�;��5��J���9�������࿼��ԤԱz�ߡW7�+�4�+�׷������9
�P��ο1��mZm�m�2�}�U�d�F>xk�}';������=3�Fǜ����0���r���{t�d. Y����٠݆qRP2	/��'�`�`$/sm�!�Ⱥ�7���oouw�%�_��o�jY,Q���`
�w�;Ӎ�\�$�t�JtP}_y��f��lyd��5�޻
�AT�%��p;�Z�5�������Jʪ�cY�k����=�v����2�@5���X�0���%B=���SL�9��UVHG>���1f!��ܫ�T�{����=����3����J%!hw�2�o�x�,Q��1w��%�r-եl�8�'��RƦ�0,����J:.��8^��w�m�H��!�b�����p�0��̩Z���/R����5�S6ń���x�qx$��T��F͂�E�눜�De�Iݬ�g�_���]'�C)g�E���K)�@�6��[�ɾl�G��;����f/�?�c�UF�S��=�\5�e���EXy�1#N?��T��&lY���(�j�R�g���m�@?���%t/d���y0NH�b�GYXl�!��;������<e�-����0e���l��O�r7Ow/��w�ԉ.L���O|���m��-�KiC�;��O���d�Gko�  @ IDATB2�qV�{�-��9�ù^��B�N�8�����u?���_?^�I���`���A��r�p�{7W��G7�.��W��z����|��o>�K�G�_L[����FM�I[�����9eL=曜���D[=K	^�┧ӿ��-jMl+\�Ky���Ȍ���,�'���ڵ�_�[���buO��������n�u�z�MjXz���qg�E/u<㓓MW=�z�^�ԉ�ǳ�Oyj�!�t2�~���C��\A�*�����'�O����WágP�t�)`)�������Fp�V�4��y�0#�)`���R�=H!���-U��i`�^h���p^r��F���o���e�ӄB�Y���$��b{��|�nM/����H�#��go��YA�T6���m�ɣ���K���S<�䷿�}>6���F�?tR'�½���Ӹg��hp�]����������a�[q3q9C���=^��/���)��i��=�^�Ɨ�Y��5��ȷt?�m&*�Uv�햾i�w��?F�q���;�x�{-���`�@c�w�veM=�S�2��.ޕ�	���*���/�$�z�w`9>I�H�-������������-]��4?�s�un�
���`�=��Ufn3{�`����Ƌ�6��t�{<(n�8�_�(�����d��t�����i[W��^����p�aڥ��-n#�K�qg��o}xK��f�9^�<:g���J{|g�̖�	%��Kg��?��=�e�����5�+f~+�^��#�h��r|���?�M������q�B`�|F�S��~�ᩮ/�O��|�k���L?��P s�ckU���2*� O�Q��xj˄+_�y���ِ����4|3������i��Li��^)/�Z���C��D�יp��t�ѥ,$����柋^��FW$�ݼ�� ۺ�=�s��K��y����t���h��ގ7aXn��L��� n�,��,�X���'�̽�&�|����;t�غ�.l1��2^����y8r�h�;�n6�}��?��S[`Z)4n2R���,���K�U����bUS:��"�B)��e5���ҥ��Bw
����&���B��t�����j�T��u&��!�z�ï2/}a-W��^�Q���D�~�`YK
R�r���ɂ���C|������"��jQ��c=Ff�ʰ>����[o���_�6[�>��ʱi���Ra�4<Y
w����Ը���w.1t��3�=#̞� ��Hg�����ޯ�K���J/γ���囸�N�v�ע��[���qd���V�m���{�g���)��l|�-t�G��,=���/��y�v+����;� �:O����1�J>9�y&xP�*��6r`S�Ƒ��ݶ$����&v.� %�h���v�M����ӄ�Y��M��[pdZ�u��c�t��.�Ѡ��������]I�$��h�%>��&�t�����ܚi��c>��sW?f���e���Om%�p�W�-ފ�^��N�l�J��h���-li��Uxa��H��I��l�J���gi �Ӝ��q���kx��&�`���8���s���N}��&ײ������o#���M���'��C��`��s��?����v�xś��S״�ˎ�ORH��n��f���wѧN��Oq�bpMW�:��g�;���l������-������3^��\�a�ʍ{����Yt�p?v�2��z>2$�۰�^�E�mp�G��R)z�K;y5�|���|��<պ��,6�ˣf;^���7^���v��|@X�Г7������X���6ڱ��~vs�����Y={���1��q�l�����i���(m8v��`��s��߻������a����ǃ�G\�0g�������,��j3�l>��oO�����^ߞ���
���+���
��`F�]��Ӎle+�6VAg5��)����&��k��x�?�x��7�Q�šI6��+;8���yY�#in���g',	ofհ<�g�Ö)��[�J����Ra��[�5�������a⣟��-tx�+��s�w&^x�çy�����.���Ń=��l�4K�0#���tY��kM&N��e��=y���b��	�d�ҭ`�^���ޯ�S^{Xq�>��,̞�o7 ��y�y0uς�&�i����ta���O����˗ְٵ?n����\���˛�����#>������X�ǣt�iOқ3�P[���ol����|o�Ya�P����}����x`��#72�{x'�r�q`���ʻ4�S�MӭF�1W��7���+n�Y�����mɷ��o���K��f��\�ˬ#\"�)M�j��Ǟ�xn�Jc��%�7m[��l�_��qς;�F��ly�l��-?��?���h�x}�{��M]�W:(����&�p���OU�Xy䷼Vڒ��
[H������؞�i7���-NA��D�]ڪ1[~�[���lߑ+Ot���R�Z��~�rOX�^\��Q��J�=7����/���]�k:���Ml,z�����_�~�~޿�N�ik��EG{y)8�uaG�k��}��v�����f^��A������l۾�v49��FOr(�s��W�7��7��O_|�����2�ɡ5��e;������_�������U��f)[����.��O�ڝ�8�4����сz{;5~���s=���{ώ��uߴ=q�����o����ٶ��F�m�m�w(r3��A�6�Y�oN��|�ր�[%�,nUl�`5`ڈD�T��I�V9��a+Q��3X��>?�+�Ӱ�S�T.��ܫ<�������kG����ת���po�P{��P��ёP��1��j��Z)N(��e�<:ﵿXE]�#�f5$2�Y�A�Ӯ�hDL���x���;��j��~�Ӝ>���Y��u��#V�Km��d���K�i�c�F��ì}�Kւ�q�n�8+�^�z�֞�fa���[�}�8c��Y�E�x�)L�0�k��	vE�+l��x|����ʰ�s?�>zL�IY���x���SG���Io����f����UG�j��i�IY��OY|����*_|�\���rn��dX�Ѥ�i O?gç�u�r���Y�,'���'��'4�<�8����h��ڠ���%_X�49���$0B)�������{6�*�Ȓp�&n�R�����c���C����=v�2.�+�JZ;������3��[����|}j����4�ҭ,��N����,\}�Ϻ'�79�)�Wܣ>�]���3}R���S������~b��ONO�i�M�Vޛ�҇+��Ow��^��s�wX_���d�|�-����TQY|�t�!\y�̓}~f��&ph+}/�V�Ud7������,��@9���5����^z�آ��������I/���L�q/�/��H�9T���8^�c	֕!������r�oG���/�>�����η�n�²��.f��\�ֶ�_|9�=�ȵ����y�-���}������$�e�(�Ͼ8܊�Ӟ�ϱU�5vq���-��rwv<�;rJ4��ƅ�@�'��k4�٨r�f���+l[�����<��V|��2S���?���Yy�<�S�&7�N�B��?E�O��v�Z��s
�U�yȉ%�Lap*k�L����	�V�Ә�q���C1/���h ���C{k��h��(�]������Y���+�
�f5N�mс�JA�^bO=}4�&b�4C{�S�@9���=��/����Տ��9�Q��ĝ��-��Q��h;WX���4�<���G�h�?A,ZՍ�{��>˕��ʱ�_W��8������?~O��pzE�x�e�}y���K����wM����ҧ@���/?�K��k;�iV���C�k�m d��M:�|�j�3fª�*��^���f���-b�����K���O��^��gW~��a{��Y'z�-�����%n߹��/��o��O"���i��$u���r�:n�T.�#�}��7>>��%��wp�4� �?t6܉�~>��_����w�w�����[�O�����FO�,�Y����$n�܎�;V��t:ɋ:�^C'a6�&W:�t3���Y�`)�Aւ?��V&������J/镍O=��(l�!�)1F�c���C���64�s\ b���B�4t�2�ǡ1|6�V����M߫�K�3�I�Q���g��ߤ%F�"��7�0����_݄+w���O6��<�@WX�I_�x>����c�`�sd�Ĺ�Gp��zg�0/'���/棱��n���{�p#�D���E��΄mѶ\]�ӈs�0R��dx��4[�!�� ���h?��/��\��[.fB��/�c������q�?���"���U3����З��>�-̯m�?�q��i���A{����w�a�?f[�ѼسXv��g��ϸuj������hW�
��1��ṗO���Wy�)��Fx���,����r��3�^!<�	���k*G��q�����TD0��Wi5�6�H�� ��1��x�ڼ'aϪs��b-��#�/Ҥ�S�>�x�)�U���I��4���Ǵ�~~��D_��L�Gw���!O:�N|�I���w�c�4�X�o6O�Z^�=��%/n]'6���p�q�u��ɐ;G�}ze;�Cx�+���(N}�g���-����ǲ��Ŧ�كn���/�������@�v/�	s�Ib���.MG����>����ǟ|��>���|�Ŗ�U?��l�}����ɣ�+��N�k�}��p��Y��i�'�*���Q'�~`C�Lx����B^q��A�/�� �A��Ξ��?����7k���n�f �L�;�p�|�����_y���r�a����Y[��Ğ~.���x��	(w���v}b���K��6�Ǿ{:+��K�-���=�qK�=��q���<�6�q�����WK�����a��t�m��׫i���?q v�ӂ<���D�W��[�}O��N��ؑ��B�K��Ӆ�X���I�<Цl}In�n�ʸ9u�}M|n���L���͟R@Fz(O��R|ӤO_G}�o��;��{.O$�U'��ë㈩��ׇ%�צ�v�a����	׉wy|����S
۟��>'��[��®�ɇQɥ,����VXhy%�箭����f��x!Ce��[�g��E�7��67'5ť��3C� i��=ҲF����Cd�2��p���'?�ǞK�!��l�7�p���S�m����@V�7mQ��_p���>��<)�}�7S�.��Z�]�������7�s�LZ���L��|q�u)0
5�i�r~���'ݞ�J���}�CߟJ2��?���S�ԃ���Cs����b�Le.ߑ=r�?g�c�IK�aj��0�v��<O��J!+	>&s�#sp��v��9�����h��א�g����֙<ܾ}��^>(^�x)���l��h��t�g��o�b���ɝ����j�G��M��Qڥ�n��7N'�������������`K.���`@��-W�:� ,YNipN���_�����Rz���7[�7�u�7n�H��?�����)g��������t�0��/-eͤŊ�x���URV[�#w�ͳ��6}Ŭܳn�m|ɳ��*�S�v-�� 1S|;G6,66�g�
��Ui9״�6����(��
�ˆ�gݞ^��+>y����,K��l��/�i�F���v�3̊3���ǳ|�������ђi���ŵP3m���M1=��`��}�ȳ}������=Li,�iy��g��u����|�LD��L�3p�e��U�ʷ�V[��2��u�d���¹�ӧtr�W���i��r*��ү��S_�0�a>4J�o��,�y�/� ��n�q�9����ō6�:�@���@�ڪ�c|ף�OEK��9tׯ_�Ӛ|a������X��GY�_[FM>α[����ʠ�v�+�_��a޹x�	ţ,ܜ��#	��ù�����_�><y%���y��~��/�r
��ܟ����+~����^��������:�e2ñ��X���Qk���d���P���1��|���xLWW������y���p���?�غ���������B�J�$/�D��G�}�#�)҅����O��
��c6+���=��~��a��T���+`�8gS[QA�6�+�$h\�3tYo*��'����w�I�2���S���<2���Jj�����َ���s�/]�R��d"��~�_�"�e>lf��>�;+��~��s4�����d�ͣȣs�EVU<�<������bk���}��������Gn�������>���i覑L^{\;��d�Z��z�W&b�!��ɢ9�6���9ǛMנq{�>#�ǁO��E�����Bc�ΙB'�
=��y���ن�r�l����U��������Y:M����εu��6�V�rы#��SW�+- h�t�>^�UP���ڣ<P�t��s-��M°���rên��G\6��С�ֹ�Lx�V����wqBE}Ov�	l��{��n�+��������~�μ�;�	�~��}�����O�H�e�9V>>�����!W>�������R���wJ�V�����9�����W7��Z���;	�S��r���`8�k8�=���A�\�G�'��4%s����^���ȍm'L�8��؟ܡ���nePa�M���)J�]a>P�^\Z�Ȳ�)�6>x���9�)0���N9�e�����V4�-״�#n���8�՟M�AZ"�x\����gi/%z�O[�#S��oRg�|⭅�]����Ů��������$�e �v��������C�,���f`��`mp^bZ�.�|�Ee�M"�Ym��;ܛ�kU֗�[�9��8a2Zޏ��*9	h�O}b����ٓ��{�LAo��E+����t&ò�d��X��{p���:������a��\�B]�vf�1��{�����& �=��{'��s�ԷO�j_�/E&��l���}Y�m��Nno���GmS�G�5^�����"e1���<��ݜ���7�x���[�E�G�/�z~�/w�VZh���������7c���q��,(���q����aՆM�r��0ߠ�d$s�ԁUO.]���RrT���Sa���a��m�G�,<`��dB���Ŵ����|]\Y��ܿ�q�|%;�'d�z�����{f�3���H�*�����[��毗�}��.�9�E�2m����ٗ�]�<y�\.<�k`�^�<�l�ʁ�Sݝ پs�Xm�j�ccMU�@��2V��ᤍb�o��R2n5F+��O�1C����wF��ػ6:�������[r��7���u���$^�u=�|���ʰ/إ)��������Yr=]��`��BG���Ӷ�:��l�2̤��I��6��Ք�>�9����`�5y�f*��b�#l����;yV��K��и����Q��ؕ�4��<��H����#g��Hwx���&һ������:�����}^U>x�%��_zM߇��.��EOkpT�i�5EJ�t��Q�S���K�O�G������\�kX�7�4g��{4��|��o��H��/�>N�-]Ǥ3��η&�{�{�k��[:�I�+]���^MF��s��9��W�B�x�!��ig�g��e�$��k�t��r_y����?��c���,���Z9z/M\a��M;+\x��r��uF� �?�����r��7>"�s�+�)�t�����;��T�n�,^���W�NN���l'�V>̖��+��ɏ���d*������sǧ��MLfp��VB7#��y��leS+t���?in������:�ق˭:��ӹz������8�ڜ?��{s�a��������������|�6#��C�_��೏�� 9t{]�v5ǳ�5O�_}�F�2�Hka��lM�t�V�|��B>&�G��fʢ�z�}���G=7�sp�x>����(�r�IN��/-�6���A;�t��,'�%}�ʳ�wi��k+6%��<JK\��/��ݧ�A��NZq�������Ocy����T��v�Ƚ�-�?�|�V�U(Wc���_�fj�K�g&|��+��
:^s�r#��&���v�VU�#�}�5h:5vȀ�ʣ������@�3	�����e�1�O]y���/��	�/���r�QQ�du�
���*ih�wJ�d[r2	��-�>���c�2�0��h��o�Mr���3��zmq'z��#����.܈p�Qx���\_'���
CN�(�.�,�w?t6�4�W���Y�� ��M�eǕVM�0d��YY��+�g���0�����a�/���O�=Lg��n24��_�	����O?��k�(�3G#�,-�Ǣ�!/?O�2!Y�A�Jl&�i����=�=�ƍ�b�Q�+"ț��5�i;���Ǐ�}�p��[�1�V&�?�6�L&�:�Z�C�nKs�g5���r��)F��D���ĝ���z4��[�����	����1����VW�{��IG�E:��L6�vt�O_�$QّK���j#��J����/�����������쁚��;�aC�;�V)vXu�@��0�6���o�^�����':K/⍽�n���54�O�)����X�3D��eO��ފ��	w�3k1���d�-Ja`�̍�o�꯾?�-z�ŗ� ��w��lޱ�f���j4�8x���/I�Ap��(N����|���^�ô	�����7s��O��l%΂�N���v�tNqk0���+�W3�z�W�{�ռGq�p����v��S���ݽ�'�}<<{�'�iߟ�O�&'��?�� .��r0��+x�KY��'��I���H�C�U��X�X:)[�r{=�廴^l=�.q���~.0l��$��8�Z���+�+�	�g��pWK�? ����@��J|�P4����/=���Z�mTUI�d����`21C欌�����O98Z��`�__�4�^p��k*�Vy��44�G{s��ؕ�j���-��Cc�G�>'�/�q�v��P'nO{�I�=��[Iv�j�|I|����u��thV��Z�_y`��7�_�T��9jP9��By�l5��"�g�>an�>/�s��j�1oW#�}�26+���44��>~"�S�����iϊ_2~{:O��N�rz�b�e���n�#�TsTi������4�Ъ$"�Bpr8?���ip���M������&&�P�n�5_mM�>�4}��nV
�d�ץ<W����c���>���&G����MS?��U����&��Ӵ�W���O���\�Y��
��أ��Ub7��g�����&n.jy
��S��Ύ�>~O�h����.n�>�o�b���K��Н:�2���r��Y����K���,���f�gc��Jw���*���oc&I/�Qs�C�p̈́ q&P�L��44VG'>M�HG��dK?
���~]Of�����Nx����^�k�/������������5�x��+��/|u��Sn�K����M�.�\����^�Ѹ���9.�x�fd�}�|!�&}}���/����S<�^
:���Cg̷���d:����K9��;w��ݶ�����~tm��7�l���U�q@�e8Y��đP�7����|��id3�����`c�.�ʘS��:��L��G����>/�7��x_��.z�����D�ghm~��=:����`�s��h>�ֲ�ۺ|��T(Z�\��c��B/� �K�W���\�L|��
�?u�[�U��k�>n����)�'�ڣr����cзo��?���ɮ#���m����$@�r�;ݐ�k"^�x핮�7��f8�ނ$KxӍvo�V�:���8��T�>U�*+3+�e��zQ`�t�wE������p@˫3� tf�����9<`�1�8|��Ȕ�4���aj�R2�[rq��n�x
]5�|�,�b��0��2bO�A��ں�YV����a";�w�{d��:��t���y�w��I;-l�	Ǟ4	ÿ���Cy�~}X_���	\�{�6����7�#�c8߀��!���{��؉�w�^Y��`�ܸq�ejJ3a�-p��6��p~���T'����g������e]�L��A�AA#�I�$�yH�/����a�k�G�I��i��qY voz^p����m1���_��0�*�#��>ƅ�io�jp��L�.�?�7 F���x;;�#<d����p&&�!t��+�lF��]x�v�/��N\�yEo�s���{��p�(�ő�ɓ�#,�g�!�����=)nJ 
_�i�E���΀;~�
�#3μ/Q���4�U/�gwKNM�x��C�ǒ/[{~���?�ŷ��{�:Y����f	,$�{�h`32���nu��^bh�bz�ıtH�GmԂnMz��c��~�[}��\�I��N�ab�؄a��C�S%_����;ڴ۷�`E[�n7|fbъ>��n>�#�x�9:d��]}���D_�Ѿ&���#Q�=o��Y����X�9��@[f��*+"�a5���c�sM+�e�,s���+��3���;�5<c'��� �9c;�Y�!���8�<����}���%�\Sw�n��Ĝ2:���h���ӛ�V���0ŕ���̠�ʵ�8����1�__�H
��_䲡P��T�>~�À�)��d:���M8��$���Ɂ�I���b�^��� Bg�/q� �
���H���(t���멃�j8�+%u�]�@�G�4�(��w�DBӼw��Q7���%�^\+�O�!J{W�����t���)Ep\6�*/|�+>~1�*��O��O�c'O�N�8�	�����;v���ZTd\N�t*F���P:�F��0�]o_�k^�<tRp�Y�[V��L��X���%en�������ܢ���Yp�+^�K\�1�P���������:�`>��<%<������ćҽ��/vP�ؖ���bR���@��Ѳ��@8\0�8�'�*��7��>M �ބ���w�W��$\�3p���+�������|@�'x+-� �ԑ�B�m51�C�,L�N�4!�D�wm���c�����n�6���~��JO�����|Z%��D^��������\�l�Rk��#pZqs�0���8n���s��i�D)�2���������Ҹ��j����
Ŗ���h�-�~�O�V@��8� &qb�S?3��	\n�>f�9���F�������j�\sa
�O�1��zậ��}vE�� �k��[�}��m"8�����_�v��G%U�3�Hߟ��6[���[?��c��֐*)p�ȆwO=��J,n����N���yGʁ�m���@S,YCXx�}/��J{G��~p�L���1��o�z@ޘ���iy��d|�YA���}1$x{|��L�����U�/^���_�_��G�,�q��_?���#7�m��/\U��.��ރ#�yǘvk�Fﭰ��	��3|P��dM8�"V���V�L��q�"n�'7����AEL#Je�7hV��|`\ʹf1��\ۙJ(�
<$�R�r)E|�Xn˻R�hD^��ա@p3x������Kd�?�CޝG ��0�1�����O]�aq�c���\{�r�ݰ�B�=��Ln�3�${L����LXl�0^n����+��`3ߍ4�~�N��{�;v������zT��ͺ}fA_g�za�k3��@W�?�w�֓#�zB�s\�xklN�i) ���
�;[�A>����P�ջ:��A��ޚ[�=�ڏ��0�b�����D���i	U�)W	c�N�����?��&���/��eOKEE <��qz^PO�m���)�e8�~�������^����!��1���n��
��oV$�mqa��YA�<YQxi
�l�����<���	/.S�`�	�__�c����9B�=��#���x�����!0��9��)�2-�S����:�Qg�HF�f�;�n�Y�^��V��z�@�ޚ�:�����%Yh%�[�����g��?��Ұcς��s��?>T��ɧ��W�n[+}��32��i���2%~�?L��;uۜ��C�򙾕��/��}a��\���	�x��\�+m����p���D�6���˚�T^f�2S4��H�A�0��J���(7F�,�A�7�Ơ�oR���WP4�C�7ŕ�%����0<'�������e��橛�j%�0��?n�{c�����c���`"���.�����1y�>��n����M�3iߋ �-+F���ȧ9��������$~1]��F�IH5���,�n)�)`��؉�w�j�����>
>4��_�R�7���7�G~��
O�3KrҰA��E�qU�_"�������+�4l��2W�mR#d�n�>d'7������{E3~�E�:=����;5c�}��Ä�!�=r���r�0�e@��VW���;�1̠�owkTH�)�m��`y�8`�5+�._��8�~�<_�Z&�%��c�!��ph�čݒ�/�A`��4�v�,wm`�H�ϥ?8�'��,��Ŭ��[��;�$��vv�q��ql]آV3h��y>x�^�4�|��oX̪��L�4�(}�2o�#��`Bv]�;�u�IXp$-	��l�cpWܽ�R ���qGA���$]õ<LX�	��_�b��GXw&�8�v��?��;�d\`�<L��ځ2eG����8�������������%͓�k�TNcz�&~�NȨ`<$Mr�'������*J�(_<��T�O+��cV���y������so\�\׮�ns�*������O�_��W��g|�QV&����kIm�|DV�-��՚X|�A���7��> �.���6�ZF]x�/�,'�Oi3.]�4���å�W��,��m^/�\���Ǐ��3^&��i�fu��ߜ�{��N͌��D�࡝��B�l��
����Y=رs�pP�*�I3r �������~D�lm��I������l����q�^�F����	� ��oD��2NO�<f2�����3闸���~����?	薧����g2�BP�)���,`L�����gY�u�X�UktJ�?�`�0�i�b�/V���DY��R�h���{e`Z��s@�{�eª;��5�6�jL_��*�/H��35�~N5�m�`�
�mM�{�Ŕ�V��@�K�<��$��̲v�e��۷�ƈ}Î]�G�c��9�+1��K�W�,�Q�Cr�Wfk�6�Mkfz�=s��<xԊ��Q�=x��#ˬYqPwc��k8�@ 3�;v�
%{C�� >f�~���=vҍh�q��������l�=<�I��������+���]ӗ�/�v +���8��t8�,_<����5�-W���l���	Ou�}��MY#=�_Fnɔ0��!���E�3 vM�3/*0�����.ϩ�"~ά�&{�I��7��<
W�)�f�<H5ʅ@���^�2oUnG���7��,����ʳ���)m?q�0�V|���Ъ��������͛\�{*��;s����iZw��n�i�aimI�V:�����Z�h+|�8	ud��'�Z����ȎmX�
�Β=߳�;3�΁K�?e�VI�eҪtJ>�~��B��=m!|d��
�:�Vc��iW:�r�ސW�����Щ��P��TT�X�l���1oЊ�=�٩yV �A�+��/q��	2��E	>\H����4bȋ�
[��?7��N�|!]�g�8��je��M�܉y��	�����y'O�r��s��⇺��G.^1�f�����8�&���6%��� +F^z�P�Dk$�F߫c�K�iB��e�8��S�ς�7Ê����p�)8ʲ��8�7Y{�(�)�I,p#c��@_ )ې@�ƥ(�L��p����%ky���ʯ�5Y�dJ>�����&�(_TN��>èvm����ogNd|i�F�nD5Dh�PvHu���h�������'><�V@�.kȾɠ�[��zq��6�p�K�Umۚ�-A���
?q��]�w�,/�3ѱuA���94��߬�n�\]�3�]�!��|m+�Wզц���̓v���Mf�罊�u�t
*�d�y^�F�Ȅ�{�cX�l~�.�v�[K�޻ś�H>��w%V�;�W-���_�c���D���S�{_��A�ڂ��;��/����i!��N�5ߊ*���r��,S� ��N���(rc����Q$[�A��'�ҝj��K9�I?�nV���	qh7���~��R6i�Yy�� Ϥ!�q�<ō	|�'����"c��Ǎ����5߬1��{�Bu�`���Ȕ0��H���I��GC ���t#Z��8jh�Jx�����X��]��ܺ��4s�����&>ܽ\ƅ^���J������@���:;���8CBCZ2=2�8�VY�C���WC��|;�O����3l�M�k̮TC=i;-� ��V'��pc�N�Uf�����G;wm�GG~���#�Ͻ+�����4�4F(�w�Q��}��u�� �6IN�I�A1YC���^A��@'�o������MQf�pT�Q���H��Қ�x!,�R��?�K����?EWT�g5���x�@�>a�Cd�C�6u�1*�	�y`�L�u3
��zE�#��0(���cXVآ&�E�+l�z��kQۘ��V[ڠ�lk�>uܤ�2ZF&����z�V�U)@1�w�~T(w���,����,���;L�K��Dj锣�K�û�=+Ίv�k@Y�a�O¨�t����`ԗ;�i$������}��<�U�3OM^&��БR��"K�~%�!BPl�_�%�`�kI�d-�M�zS���.�v�7��w�/��BB��.K\��P�+�*+-T%���#����0�*e7(i�W�L�2�����W�M1Y�e��=}�}`	�X.�Uϴ'��߼�����÷b�����7x˧
�LK �3���O<���aKS� O9�mDC������/���cj�t���q}5���r��z?�Yi��2�|��Y�+�m��,מv����VmH�;�ؔ�&��~jj�:�,��96�ۛ�:����D�ѷ�Ăei�LH��
��u��#r�=�u�����՚У>q���m�Fʄ��-o^b�G��q���=[��8�ҷJ��B>@�!�ԗ��:�}�b5ʃ�p�d}�
.���=�>y���=|*=��'y�������P����8���9�����cR��$�a���0^�P���\�;,�����O���{ڦ�NE
�Й�5Ӻ���2�0Tp��'� !���yo��NM�1�A7HG����ެFg��]�A�RnT.���
I��F�X��Ɨ��Z	�ᇇ���p�JVܱG��G	�h�H�@������/ ��_K�&�
�l��ߺ�􊾃��D�<�e�p��Qm�ڣ|�T��M�!#��L
�~(�iV�N��e���~�8����Q�l�D��I��;�|�w���(�]&��c�뎠�e�K�=XP����=�(�Gr��Bċ����X��_e�����q��Y#"�GV����Ҋ�lԻ�@�Nʞ�5mĆG�Sr����]�H9��{�@Pq\no�ns��:L�U�<�C[�*�r��l�Ѻ��@�-�	���q��%}폕2� �����(��YiѶx�d���˾UKe��_r4��yb�S��.1`�붅I	��d��<~F�T�����l�~1����`�i��⃟��@��Y�6�o������96���M%L�.�9�ʴ�*���ٶ�K(x�o�T���V�0\�GaU��¨2 2@Ϳ02�Ș�X�B�
薩y�%���V�I"�Fi���ʘ�M�����oI�x1��� C�h�K���~�W�����'��
�"ԯ���(7��o�	3J3���.r���mL��n��5���z�0H\�9��;��2���M�Ҡ;+�p���Ƶ���vIŉ"Lfu1O&  @ IDAT�p��)�59l�m~�K{c�V�f�5a�t[R��<GR�A�����Uc��"%����]]wm|�Y�.J���+̦�oN�|K�ʩ��e\�@xqE�Ԍ�W�U���{�5�������8߁�2�W_7I��֓x�a&i���wG����~�!�B��#�z��f�c�aNp�;��'���ar-m(c^�oށ5�4�ؤ�rj�.��?�:N`�ݻy'^���	��4����V>�~�o�r	 �>ߒ`&�g�{(B�G�g��R�����{22�4d؁I��&ld�<��Ue��O<�=^2�͚IX��Aq50l9B��
��B?n�X����}�ު U�3+�I�z�*1�4$�ei�ڇ�e}e��熥q��d6��t�42��Ռ��ۋڿ^_	���d�~\9�������m�W�̐�.�ŮA
��Q"������xhi@1���)\���,�bH�|2t��-?4��O�����.�~q7az<''<a��⸱�>���	�xx�;6����Z�!mո'iC�5�D܆���V��AP�-�woHi��@�=�����3� ����ߓ��!�^�х��`$	�i���ܫ\��	�eU�]/W��Qr[���8h͡�)=+3�J����ɝ����[��紙��J\�c���/\�bP�
ޭ(Vg�JŴ|Gx�7���r�rM,.J9Z�x)�vk��'�<�����3JE����Y�K�'x1�����<V�#��-��r�	,��F�(��>�|�^}ޘ��.�o���7����1o�*o���ͪ-Ő:I������x!�o�A�"M�ڣN��~�/�	�֐�كJфw�0yR��H���C��%�d���y�U�G��`�C�Et��ؘ�;�Յ��.�'^����O���G�yK8�a&i��Y���y��8�2�PVi��=�㤒�
}�\e	�z�|%��>�r�T�V�'�@��\"��
lx�rJ��t���G���߂��	_ "|�uZ?}2m��F�� ��S�%���lY���p��L��>�/�*V����=<�عs��1�o�*<q�/�@���ZFVz�<�hR�����Ʒ��<n�"�]���x�\}<��Z`^�^�<�v�R��˄��ǅ�`��׬��?B<zG&�e>is�+�<����yJ8<��;�� ������Yz���_����<��gW���I!�6(���ڜ0��7�&�e
��(���?L�S��N�?! ���+�x&�w��Y�[ܬgN{'�݄�Ee�sP���4�\G*{uBY�g�ԁ+�q�K���#�'#�-O�6O����6>�ݸqsx�w�m[w�aXݮ'^/�iGo������B���93��"8ؚ��~Ka#��@4��?q�9+��7�04��~���^�*�7�,-#t�`��Qq�m^���5ڍL��Ɔ41R�jF�Xip	)�_*��TN7��FaXa�n�t��g(�d�N�(�ap��
kn�
�O|��Jo�a�l/�(�B]��|]o:��JH>�/*�NҀ�5)
%-�W2�?�f���NwUw�;�LK�
�Y�9�R���s`����2C���*O�1ɥ���Q�s�p���/د�2��:+'��G�Cm�D"��>��@�/q�.[i���Gi�z��L>��'�P2����Ց<G���6�	-2�)z�F�(=xS�M=1��6M���x�C1�A���� #��}G��N{�0�Ey'���8h���Yx3�KD��&F����Z��58�1y�a�:�&���5;�C4�kU�<��]��l/�>��N>mS��T��0��s����C$��;&��KX��?��?Op������3Z��W��!��n���w�S=h��C�e�b�)��^�r:<P-.�S�Ȼ�G��>s��_K���#��8�mN��+��3�2Y����*�p���@��la��h�3j��U"N�<�k�Q���ċ�_�,���wo�R9�ä�x␉�-����f���8����1�o1R\`HÜ���i����8v���+���U`�#p�us(`�y�U��"��V�-ܚd�"g�0Y�"��|���C�����Ȏ���cf\�o�U$@>�X�]�|1(Ȱdv�{�/��U¾,�M�Z��F�XH��x��p�������ysZ>_�'�ӠªaQ%�7W�q��k�X�d[�5��e��Nl<��ʠ5@ZPTc���$Q�nk{ȕ+W��q�yǎ
S��g7FL�cb޻Y���Ťa���߼�۝��1s��[�����۷�Liݩl�Jy�I!&�_d�çaުe^S:��;w��/]�<����'�|b8hH�	��+�0$B�����T�~uf�Ǵp�Νt����A��`��)*��/7�y6�ɍx��r��%�t�C��T�b\�F) ���/��kh�~Tf�O��Ï��t���J�*���|⥢_�F˽��O\`���oY�_�
��]c��d��:tK��>���h花��Q�"��P��,�]���y3ަ8&��Mzb�x1�AI@���jC8��8�O�_˛|-���µJ�����L��=�n�~Hy܊22�Z�����7��x0�e��Va=�a����P\�>�)��`N�<��3���1���rQ��@݆ghd8Ћ���,���m�	��� ?��E�h�����i���Jg�dFx��XƝ��x�u�t�_��l��ý�m)
x�Ͳ�<�����c��81��ҁ	.���B\�x�M�N�b�|u�)*�ҿ1P�x�`���n0�/@��#������6rft��,^+Ϡ�k@������I�c ��-�ޒ࡙|v:�b�t3UaU��%� P�x�n�7��W�����O��e�,,k��	�y�Z8|��Vlׇ�W.����Ixg�ߨ���ǒ��I`8�a�}�d�<$<�U��n� #d�;-�g�)g��E�g$Wrj�_�'~���YF��#<�β�%t�o�c�wB&haqc���!�����߷�	 �>��N�����ܺ�i�qA���Þ�������@���qE��1�)t�1Nbv����:���5RjO�[8���9u����;U �Flre�B�Ki��Q�5�(��^��̺�_�f����S�=��@��mO��z~�6���3Bc�M��������+W�i�В���(x#>����:�|^�MguFp<���:�F�$�+���NA�?���|�xЈ�̤Z�GN�ۦ�+�Jm�;q�Ff;i�H�Jk��/�������騣�X�dK����NO��t��鎖��DA���������1#��?�d��Ӑ^*�e�͋���!���C�ˋĘ��'<� ���fO~��Q��?��h�>7����I')�>���QU���in�x*�$2�����ݿ3�	mh���/�qz$ޖ�n�s���k���kP�|����\~�b��l���/�zg+��J0��D��V�Z��$�e�p����9L��E}��`�r!^�q�f�Z2�f�)��H�M�#m ¦��"J��m+J����W݆W�^ɀ��D�%igUxߕ��{���8"K`�Ǆ����%���(���]kÓn����ɼ �NN&`"U�����W�|�Ä��c'w>���7��G�@ܱx��~`p�8�]����#+�����_k/�Lk�I+��k�O�C�Gʔ�^���z�/����S7ȥ�Ï���u��*�|�mN�,h%�q��y���%7��`[	��%`���� �hm���@��5<����-�����,�h�#�w�
���)+Å����+�9����N��c��֨��A�:a���;�=�_�O�q���ɔ\�S��� �C۰
_�g�S��y��x"_�p�5�
�`�`ekYL��_p�'���ǎ�`��'�c����K��p�<;�Z�0l�w�
�����L��dU�q�L���㎁8��$(��0�ƥ�MM���q����u0ЭʛJ)�I
338����aˇ*mnY0j�������Л�PV�G�<Wѱw��⬪#޻o����顇�h���5�
/l^�9���?��4`Tn4��Cg�;a�O}��&��	pc3K��Spz,�<=�ʇZ�fe���������sh�С#�N�ȃ����g��zl�):�7��t``h�I�"�|#7�Ф�n۲lLh�]~������U�ӡ`2��;�sړ[|H����4����`�r�W��=��1���n�i���+��~�LG�|oF:�'�^���<�;*}��fMg$�I\�2�,����KW,*��o�T��aǶ���@��T4��&��fn�cv٤q~d�Y+l���;[�z����z)�HY�z�,~�
�2�Y<��N����K�!�!���l��#
��Wz�^�� ��l�|�#��挅��fW�x�/e,�v!Uz�y�,#Ǎ�CV���rhz�?pZ��'e���/ˡ
s��/
�6���W��dC:��iw����I�5
_!��YU{��
�
E���=��L�TU��i�$�e�<pe
��F��<<9o���R����`{eM��O�Py������w�z���&��أp�1�G�1���L�d�#����E�?8�����W^� �z3͖�WpL��|��:��R$S�L�Bh���S|�ň�W�2�3���>�VЙ4K����ޱ�sN_KC�@�g�]sښ��/'ƣ4����>sfv���D��9֞�\mٴV�IiI����]��˖��{LZ����|[�t\��l�ږ���x�*c���[n�_m<q�B�����>|�\��]�!r��"? �Fl��&q�p)-ayz�{�1��_�	�o}���U���vtD*�:<9��c
*���h���x�FrS��5���Z�U)N©,��z�Y}�N�=��.��j7W6�R�(��"�-�~١e�Y���h���L���zo>D���CM0k�R8u[�T}����[ʀ����������MmZ��lՄ�f�E
��U��o��`aت�-zhD����-ձR������
�4��F��,eG[Y�0��ZW�V޺}���o��ȻK����VVBP�Q�i�0i��$1�#��w7 ��X��6+�� ��YiAyF��/<���jɚ��_��mOSS��^������;Õ�Wt�����2�����!�/����P>�&/��p�X1��?i$>fU;�H�e�W?j����'N:�����@��(��6�ġ#Y�@�{��n!�r� ��HA��;wj�j��>����҇N���S��G�P�X��s ���N����C���:���jl��{³�A)���Y�]�|���w�-�>xw�^�l����,J�˛��c�@X܀����vy�G�I�{ɑ%���U�k�6;�
F�I+{jofU��j�� ׹"�۷�|l����Cy��!=f7k@_�'���F僴�<�M�[m���C�Է��o:E<(�K��	��q/Ҷ�Jh�{Р�Y9P� eǫ�)/�-¼�D<0�0��hD��_�zFu����^�Z���q�h�gq�x#o ���m�q��vK�ңF�+%ؖ�x�;��Wn��?4��x���;#��<eP~V�0����Rm��M�6�K�+�a`����Gr��!=���:ǣ��U�iZ�&e���6V٤�K�3H�L1xT+=���D��po&�|��$�ͳ.Ǹ��K���E=��zǰ:�;�6)ϒ^�S��I<}�n)s����C�ӛ�GV�������6����	��z�3�C��u&���y�;iNzyg!&<�|�{�>�^��:,��C�>�l��ƌxhe)x�n�?��Sx(U
�[�t%�,$�`��o�a�'%A�& Tn([�킃�e�;ܲ7'=�[�ԇ@��]���Q;�v���@}���̜v;�k7�ͫ���]S�o�R�1��	�G�Wa��d�J5�i��:(��蛠%919�v��G�3�{��]��Ĩo,i��+���U�g�����<���r�/,��8p�'��E�q~�����_Ǎ���7_M���|S�����7�W[M�U^���m|1�-O�)z7aM��J8
*0i�x�����2�c��/�{�R=�Y:��chwhD�"3[50ٱEJ�v&��oP%�~����u�hA�{���l�f4���`BY��Ј/-���MW������O���[�ի�U��0��*<J��7���ʕt�+2!;�G�l��q�
���y���RI�b��C\`��"�v]���j�����Z]�'a����;����?��ug9������h4%�ѡ��m��I~��"c:*� F��|�%m�����A���&���rG
*���ljr\���P�h\k�@�� �t�$ա婶����ljfkY�v�V;�!.y�|�U����Ki�dp�Wn�`�yW9�&F"6N�M?8�� ��%�Ȅ�J(KV*U~G�&���'+8�.9d{t	�w�1tJfF|��31���y�!�o���yݰ2�2����u}����}v�W�ޔb����;�J��tDo��x�_0�3�!}�w\v���u����}Ƕ���������[�| >3�4�����&+:P�d��	��x�C�t%d˅I⃇�TU�MBF�cPn1�W������b��FiN��;Z�b��O4��]F�i�4���&M�@s^��о ���$��.P��7�9��QyP��<X.���i���5D�i���U�pG6��1��ܣ�s�B���/a(-
C	�����aY��R� oc�����A���t9�9�Q~R/XT$N��O+��ڤ ��l��HZ� k��ɀb���/�Y��d��S:��PMX���#�'�c5"~����с��o��0��le���?�������=��fe�I�2	��p�����[�R�U��e���1��������V���I�E���'�:�iKh���a@�Dxc����)����&��%��.�1�&{�Kq��iO���Ʋ��	Xڇ���.'N�t�݃n�~���I���x`�8����M�}�ח@���=~Pǝ�/⦴�.4bwA'eZ)|=�F�+0�XO�#���t<54�����Q�8�P#o
;
��R�5:%%LZ����Ef��a�Ù֊�;Ku*T��� �����;��mP� x5DRЙUc�{N_�>��p�̙��g�C?J�R ����V1S!�-�~��L|a�^�x��03�̰���26q��]2_�B�e8~���P+؆+j?���p�ԇ���	W5����4���$_���V���L�L`1毭�d�+�)0�x����rԿ�1��~��VkƋ<vg"�E�9f/5�DR�S�S+ ��{@)��>�gCK������7���2�%�Dsx���{�x\�L���q�c����]�����P���[�"'�Q40(l�c���Rl��0�����l���r3�޷o���CG�GN>�m~hƎ�G�Q�e#f�H7��y�b���;�SG>��}׺�@���Ċ��7M�W��+|U�+|�dj���os��w�������O?>��#��v�H4�-+/����y�zNo���p��ᣏO����*'�2�1.'Jj��I��,�cY��f}��<�y�UY�Ү_�5�o����;��W�g��OV�Ն��jf�����e��(B�_$���u�P�ࡏ��kΥĢ��hEF�)�7�Z1r�����H�P;D=`x�������a���e��A,rfP��y��>jyE�+�k󴽭,!ZE�y�����ͻ���1���͛7�E�[�H�<n�m�k%%wn��R�s�vM���Ш�2u����܅�Ý���N��a��S�V����������ʯ�
�իWuC������<���g���b�҄��-�Zi��>�~e�Y�L��eE�L[�u��J0a�E{��w���%Τ��nx����è+��Y������7�����r�MS���G�%M��A~L��N	��ğ2�����(����M̪:v��j��O\��5�jxU%h� C����G���^�P|n�K���ږ�vX�O��v��B���� �1E�t�K��,���H�������Lhc�/��$l��8��_]�l'cVO���X�1	�w�P�2���g̯�&a:�n�&1�IE�,\�S��ԩ�'Nl����i�h�Κ�������3��K��V�A��ݹ1�H��Ni�2�@��TNp`L�����3f�G�ض]�ǵՂ
��.�ӱ�ɀ�p�>-��8a���1��/V=�5���\r3(h�������������W��7B�`���9e�fKi��4:��Z�f�,+w�����/{y���S��;�����8ȵ�1�!��i�?q�ͺ)�w��	/���m>��`���e�Δ��
�m��t�����7B��RC�¼S�R��������p���N�a8r䈯*D�O��#��uƁ��2#J�6��2r.����Î�;|�׵k�����aɺV-�l-ޝN�Ur�wp���͈�syƬ|d<��)��j��ʪ��Ķ�;����a��v%sf����ߗ��J ���=��8:<���g�}vx��W��V�6/�O-L�n��h�x����麙�e��y�V�ȟ�'��/�_�xqx��u;�{ÌV9�"L�\�q��!<�}�i�.��|����?�VE+��߲Q�c������Mzy7�d�p;�Z�Ǐ���
��@�!r�ZrCi�P{�2���md@����}L�#�Gm����W TቸlM�JB�)��|a�?�nh���Tb3�+3����/�3p۩r�����N�8�:Q�p�>�W�_�����+���ڵm;v��MJ\^��ᥗ_� �1L�#�=-
J�c�?jz��������p��m+v��ǐn��E��ܬ�0A��Ǐ����d0���������Kw�3��y�tXFZyQ�%�5�ͧ�~zx��o�������~���o����4�K��J��E�����7b`��C��-��U�#�fl�7x�1�0�m0��� >ؿ����
���8I�� ��^���+�7=��1����pld���	�I|	(���?y(۩��-���:[T�ӟ�v]�$�N�o�ւgN��#����x�RK��+��UqT̈́���
�_\��~��IQ7Gf< /�r2rD6.W���(o�M�5$�Y���K��;�^6h /��>l�	����{�x�7�><8�~�À���$�����e"��b2;n28��c�\Px��d�d֌�0�7
8�^����ܼ^/�g�U�����v��e�a�6������uK"��̤zư*�yWi��������gV(��ieE�:�ǳ��O���,U���|pǏ8�&���uޤ���eY)7^lL����j��ݔ���-@�R�9�Ɍ���G�r�����d����"���e��d4��v�%9�,66t(K�o�aO��Щx%ʊ���2�8���-����=pl@qؽk���˯i��]�Z�$������z8�����`����A��w��%3�"N�81<r����bH��曞��J�]��[�}��'��I��H� �(�(������@����=���ts�A(�/���ӧ�N(��5�y��q�=ycMWy��Qr"��l�2F�#+��c��l�C��P�R��7|��v߭:�>||���O���t��A��C�91���?y��a��=N�VZ�~�mς�ń[�Pny�MP<����	FX��ݾ�U灶�~�D�TGf�A�<�t��-h�3!�#ҁ�zCڨ��@	!�MZ�"ޢZ��eh���EI��G�s��֫���������j�*��@��U��vͪ)R��%�B��UuV0������rҦ�Nʖ$�I�g��j%�Y̶�V9�fBxV8�O���~8<��S��R�*8ceLe��V)n\�╜=����ȍ�����sU�f�[5����}�����w���wg������e�&9P֦tK_�Yi�����n����k������$�CY���㏴Jun����H��Y�D����.8�ox���5��5����W�]��������K$9=���8_������3�@�	２^����A���O��\�p��y������� .���>�T_Pe�����C��˵�i[��c�I섙W ԐǏW�mL^�����Cw��8Y[u7�H�I��	�^G>y�C����|Ȅ��1~�ӂ��|�Ւ�	ʺ��ZR@�K�b3p���R�P��ak>�������e�v��?�O��EN� ]OZӇ/ɀ�/�
,����������&?j��JfL~xrG8���0��x��"��%��{R� O���+�������Nx_I��S�)|)ȁ%\Ij?����)a���tS�yJt�<��aޕbH=���ƂWیD{F�%"Z��K�O��Vk_��HWj�:g�̀�N7i(�UIaXW���a�C�'��wA�/W�r02ue&JD
�e�!`/���#_�h01rZF�O>d;��!�V������M�q���V������wֻ�G�}��o���˸Q4��3�l�`%������~���?��msS�;�>�wA�����7�~��>���`+�P`QP.JQ�����[�R�������0<���Vt٪A ~Ω0������ɧ��l��/��8W4��5[FX�xB�?��φ'�xB�������Ib�z�����+��<�)y��Rv"���;p�?t �C^�!`1( �Ok{���;T�����r�>���;û}0��_��»����|8����gؽg�����W^^y�e���{���֞^.:`���cA�G�����u�Q���ܵC��KP�� �_,�:g��b��E�˨^�`Xt�&���`�|�3۷�����+�Fj����5���J��Sr�1�2 C�AFt�Cyc6���i�/RZT/�R�(<�Oa%�J�x�Ҁ�3�HQ�Gy��� ��iC��;��d#�~{x��\P{聇���Ǫ?�aemWӊ��3�Z�ߤ�w=|���ᣇ��{���p�Ժ�p�i8qb�d�c8$e�]
2�i��`�4�<"+�,��b5����O�Vq�V&�_�T���[`fU��5���ڶGZ���wj8�أÉ'4�\9�|�.h�T��j��͆�3F7�^N����o�������*��Ap�`������
��RᎣh���8F�ڪ��A]����/����k��bޠ7@��*�c�����cp��jg[�`dE=�N{h��7m��;p��?n���zM�=��rC|p�[��N���7&��C�c����;dc�4Ȼw��� ����*�	/��O���U�?����~ a�"{t~��C=7Ϝ�O�M��c���`�<����w&��/<�1o��ox^��o�F��������o�r	D������?~��р�� �����m`��
x�v�H
��2c��U�r��ѣ@: ����"U�7#X�s�PE/j�t�᎖�uPs��a�vUO=�(,��Z�[�i���e�Kf���q ���ו�eVx�N0��%��E�i4x������ע��*M�I�:F5�qL��+k��F���\q��՜U�Lǧ�kJ7Ե�5h0o��K��F�����7��`J�8�A-��U���� u��?�|���x�ZkQC&�'X�=���&�ѓǇ4��_�D3�'��fQ3��/���A�{�g���E���7_Wغ��<i�Ղ7u���+f����C��s����_�l�/���Ɠ�w�~K���p��~o����Ymo��S�t2�{�|�X������4Hy�{�s�����g<��裏z�����W���L׍eL�E.��ʱR0�}0�@,C��H<�N�����|��?3�˲o��\��2�u��𙶑]U��7�.�.]>��C+�|T
E����g�^hq�uh��BsNJ,[���fʛ<6<���Q���S����j{��ˢ�����<��Ӧ�;�����ТV(�x������=M�{�ˁ������fݯ�|tz����rDۨ�x�qie?�8��Ŋ/�S�I+Z�+�� 93�裏������G�Z1��+׮��;��.*Z��<����k^7�0 Y���MnN/U�G���G�%�J�)<R�q�gN
6�Y۶l��=��l;����?�a���}F��~����;��+������K�yj׮}�;m�]�Y�*�
�oUc #�\���r����?�I[JTb5P|�Wk���5�A��Xk�Ge��f�U�(������6�!�*k�����>�S[���?*�U^���"��x[[�N[$���zrx��T7#ċ���2����A�C����0BUx�`�ɮ�V)ED�L�>{v?3j�)�G��-#�f�������x[�{����0��M:1�\?ܛ��C���?���i���h���$��* +�!�|��o����0�����?�6����O<-=�Z���(�W�C�S%�.��J�z���x��߱�1]��wxO6�	#�Ɓfĳ�bw�Ý��!;�ă7�K��b�C]kM���������"�I����"�ɼ�*X>7�HAH��U��%0ԃ�$$�x�l:�~�0��G|�y�t$-,)Vc�����Spa6o֌�n�ٮ��)բ��)H��
]kɀ���M�������!+�����C�ЁGL�͋aJ	�Sᥬ%��	n�aYL5otf51|k�K.����O�jz,_䏜���4ɾ��nl���t{õ��3 �82��;�q�p�S�,��&�Z]�^��W���������D���4b��ܽ}���'����oyv�8���Wd�����r��6��믿:��?��g�uɫ�4��m%�'��g��������~�����?'N��?n\�Ԗ�c���[>p���O/�4����R���İ�ꓳ�x���j@���Z�`{�?��?��q��g?����ɓ�zP����IA��su(����IGY�2����2���n��tz��\n$h��ĵ��(�a�ef��5����nW=C�ڮ��iVX�-�ŕ�׷���a�A�耏�w�.d�w}��'�|r��O~�zd ���k�x~x��SÒwu��ߟ��s޶�w�^��@����R���Wt���-��	��|�V1�,���%�PP_|���.���4�c��f��]�R�^�@�E��iI�C�Ȁt3��ӟ^6߭!]���������ʿ,���V����>��т��m�ֽ��YNg0�U.�C7
ru� �7��%�ڪĀ
%xU�e�gE��~{��סh��tQ�%���B�� ��?=;�ֳIW�<ttؾk��Ǿr��Z!��,2�O~s��2�{�ޮ-��%��$zpFl���?^{�UU���\�ˠ~U��e��@���]��T�My��%ۤ���>L̀>�#.2� Rgf��r:�����i\�K���ѵˮ
�Je9���k}S�\�DϠ'aZ4��W�T'h��Fi"S�G��/u��W�b�[�R>�cE*���?=eb��:�m#r��	n�zw�!W�!�6&��=`�@��ɘn����>.�o�Z�^�q/�'&4������B��|Ř��G>G�r��NL�}mD�e���{º���']P�4��q<�q���h2>�1y l�&��8c��M?�����	���_�&���#����$`yvY����C���f�Ɛ�W�j�p��� 峲�~��a�K�g˥d�A� ���:|f1Y�T���)�;H}+��NVPʥ�Mm���Y��=bXV���8S���ʫJO%fYJt������ ,`Z^fH#� ��[����m���6%Y3[(_R��J��5��-u��z�aYJJ�EJ��t�T��<4ś���`&��њ�O��\�UZH�xaւ���KLd^��;�p)��yJ������<b^�%{� �WY��k~����5m{�{�Q;e܄����	�u��NjH�=��X��.���;��",Ip��t��2���(�-p*̸A
��D���{�Tc�B��%ZyY���3�\Ї�>�v���XH��1#�bF����������]����3�����n�XԶf��4(9.�SR�޸=���Ç�2] ��ݫ7������J��=�u��hx6_�!;uy�*�VeG�-q���R2�����x��������i)g+��x�8����e�[��t�����F�s�+"eK&y2i�� ;����W��H^�-F�������p)��%g���^f�}�Y+g������_�-f7��^���������_����GJ��pV+(�s����{f8����VU�ř�u�t�򹢏J.)?���l٩<��wm7�*#w���!����
�tA�@?yB����J�<\�v]{�����d��g4x���=���`���KÌ&!��F�~p������^+EUJ���Ǐ�l>��a�N�EIaE�IR�*���P�w�=�^�Rz]�Y͂�Qzo+=kڿ}���aU����^�Jה:p�4��@9�V��D����c+�o�R���e
���Vn�Y���Ђ�3���}Z�5�lmNgK���Ე�U��N*�+K���:t���=Ӂzt�i���V���aϾ��gZ]��:�}�q�:r������Xe���{��S�~/_���٥჏?Qt����<���)*&tP����:C�Gi�Y�٣-s=xd8z�A�^����s؝�J߅�������+wum��N�Uߢ��ݯ��4fi�gێ�a߃���qdx��=�d0��G��З��bC�����Qʐ'�P�fhg��︝j��`�Ꝃm�O�yÐ��	���u�s�s]��o�nAQ4�,�b�?p|�2O �-k<��(�l}�PT��,�����M������a�aE}��	��u?(��٧ 8�\�ᦿ��;
�
��>z#O*��@�<�x�E��v�oȤ�rIY�v��*n�Ӊ,�Sy���J@��N��=���I�hj[�g����������w�f�jV�f3��mP���}�S�\��!w_� �Ɨ�N%I	+j?%sZ�u�� mS*�k�9���J�`%eߡ����0��,�D^�;�	�RC�TVڐ��J{N:i����<��Uӵ8k$D�=�e�'[��'���옮bۏ�+�=m�����q��t&Wd@�K�S&���_�Č�I|����@�u.Iҕ�e�� �q��k�R�Ƣ��w(Fo��J&u�_����� ���~q��UK�
�"�(��Jpţ�#����d� r��̖1s���G�4�*�jV�9�*_����g�3����,&�pZZ��)<m���̎ʯ2��W�,{����q7>̓�7���ƿ�+n�����k9�r��g��o�y��F74�Å3t�R���{jp�vO��M��W_�B���%:�����Yf/Q$��]�la����r7['�+78A����V�ϝ�ԍ�SO=c��t@�ۇN�:�5?��O�#������}���l}��RV����SV���e������:b�Z^�#��=#~��I+@����L�S/��	������Q~(��IO�H;R�=�8q�����R� @�_Ь3�5�Ja;6<���,73�������2�k���~;��W����������9<��#l/����}��|�bUۥ3���U��_~ex�T������>Uum�;xd�W�����m�����]�R����q�  @ IDAT�Zu��w�3����߽�mG���W��i��<��s>0LZ9,�ꫯ{���o�V2hW�{�?ȉ"2���w�m�����mT�t������.]5�gu����A����}DTN�+�tJ���q�턔ǴA�a�!_)ㅧ�[�ǟ�x%YBc���?��
+5�=��W+h@���~�gVj8��޻o�����zS����Z�YY��.'�5�ۡ�3�o����(�zfx�ͷ4`X�J�9�j=���"}�}�d�x_��7/jP��g��Hu�o�lҪ�#�7����?�� �3����(�����{Q�	?U�K�$?�V2a��x&VviE��g���M������]}�>�>��d�+J�TN�38>2��H���������y`��������1�m������;��d܍p�}���&�A^��(�1����J2v󞧇� {��&op���Y��v�t����<0�'���7H�ju
��'�*���{L��Og0 uܰRz��z�:�}�'�Ќ����눴n[K�"��C�'i�"8���U3�<1�׿�?�C���^.�`��!Â����d'�z���ǜ�����J`C^I���瀢2�F���,�1�G
%�1i�\���+���Ŏ�ŃaT�)�@���dh��>��F漢*	�� �����P��c�E5�V��M���q���?ˣ5
=^O�W��c�h�=5�p�0!g��i5!�n���t�>q��>Fˇޫ��Ws'~F�g��I�a���#���>�h�D+�p9e�U�e����:�y�nn�zNסn�\nz�����k3�Z��1�U���b�����.ǒ���:QP�B;�o��Ċf�Vu�nQ��(�������S�2Cy@i��3
�F���v�Y����-V�:!g������P� ��&y7��K8��;u'����\:��n��V�PΆ��o���Çi���?���Zf��*t��u�� �=	M����oN �ǟ|B�uVۃ�4��[����+Z�|�O�yƷ���чï���Sd͹���*�!mE�(Y{����F��~o���YlC:|䈷�핲L}��m7g������ҷt>��~)����o��A��4�H��׿q���ߧێ8O���˯\�HۛN>��ˣii;3紙�*�����~=�Qۡ��W�9dş|&�Gy�A:e�
�����3�M��c[3�Ф�2�M#�(G�g�fN[Ը��ո��o��}��OR��*�	��@��Μ���-�Gy�W�����У8q����)o/h��]��j�G�vk��u��gZM�c�����>rN��W�-p�u�����O��m�{���7V$>��������	]%���e�tQ�PQ�b+��wj���ǟ��/�F+d/����=�|����׹�ݞP��*QiQ�0�d�^?�w�z�
�G�Tʪ,�ed7����Z�d?�GtG+���"���z����pp���{o߿W<�c~�[�ŏg�)k�G8�˃�y7?*�����f�Ǒ�����{?�y��3P��DMx��S'@C�����p��������2� ���@����c�de��.��/<%�8^=V��^Y�B��y��G��'��Z�}�z7<���X���x<�C?x�+V+<���..ᘤ��O��!��	8�:D�?��g_Q؞��222����ڝU@���BA#�ۉh��%M&E+����� �&=U����P���!0�G;tX��?az4��
7,�f0���vU<����+TѬ.���7���5n`F����G6vHcy�/i�M���*~��4��᪒GNE��W������<�'i�>�7�U
z��	�#��ЈLಂ�wA[&y疤������K����G��v'Wu�F��n)TG��绚9?`���!l� .	ٽ{��µl�|�W����ޥkhQ���ч[y~㍷�ֶ'N���է�z\���h�*R~R�P(���(�(`���R;H��j��}��$<2�;6~���Qޥ�|�L"�yz���*;z���҇·MgY{�����oz ��1Mj�߳o�f��>r=)J8[j�CV��_��MI�f��M��5EtiO�Hs�<7 qs�A�V��=��	��4�z����AmYB���/�r��R��X9b����&������>Aޝ�r:�-�>�}��ygp��3��b�V�9���(V�Xm�?>�wJ�Z^I�;��>�Q�5���VdrQm�&ĘY���Y�	qy�_�|�ɀ��,�	La��a�_��W�ʭ��?��������=*^YA�r��-��yY�_|���
�QT�i3Qr��a ƀ����Ŀ���?��ta�3���������A�]������C�[Ҷ���?����@�c�u�����0�����u�Aٻ���^����Zn�)���xP4~������*k{u>��_~�o.�ZU����?|��3/��V�����!ɼ�DM�igl��K4��Zސ/c@����=�	#%�^fo"0��U���c������$�mf��	�i�U��tQ6y���py��C�3�����(h�������l�{��=y����a�B���8��K����;<��.I���J�恮�A
 wz����J�Fy���;����(j�	��ൻ�#�b�������S�x�	7_����e����JHyB޸�c��t����(�B�g���A��(�B��B%�
��Q���h����i���VF�4#%<����
�h�����J�T�Q�Y������o������8�K�T�d �1���Ǝ��C#��A�xy�m�a���"w���G�y�j�U��"���Z@�6?JH5��&&^k�^�7�4h�T:̗|�1��/_�,p��Q�ь`�s�_/g{�f��a�1��/(3��ެ3�nߒb�[��8�}�K�.��V)S�n�ߖҳc����&�>c�y	��e�<�98��C��{��	���׽-��W_�+8U���P�޳͊��,�R(��ՆW�En������?f�f>�6��M� ���=6���g��U&�&rT�����|K+ lOb��?���5Vd��������1��^��[v�^���(��.ΪLK�mW-�����m��KRr�C++���1mI̊Vɝ0�k:����l��"����i��4v��i�&Y9`��_�������L3�`������ѹ��|O������8���Ԍ�Y}d����Hr5�RЉ�;�6�I'g�Rfy�
A���eL�7<��'�y�?.�:�-�rS'���dݼ~�e��Β8�8��Z]`;Ӊ�Ǉ����?�"�����J�|Jn��+�_z�%m5��߉@��9�0٣���[o{���g�n�A�i��2�E_�~��1}��_�u[���->N9��*���`o�p1H�s��2�����7�=���Jǋ/�F���i@�aɯc����;ya�n!�{؄�~ʒ��)����^ha���6<�;�NL+"��{+� y�;a؀��Lvդa�Қ�g�c���F��z
o�������=�w�?y��V��\�?Bn�����-� �!2e�+�C�WxD���)�L�`�:�'m%��U�&�ƭ�|�S99P?Y����v��ؘ�c;���<��x�.>H+~PLX�6��ǣ؆72�V]�wI<l¨o�a��<�'���x�7�!	 �ȻG���݇}������p���}��4TԪ�U���OER3dUUR �])�Q{K!(�:Lv�pr�`��P�1�@�*�� X�262 ~��h����eT7��0rꅞ̉i1�� 01E�������\I��\����~�M>#�$Xf��n}L-���癰�E�7�38��N���2�;�٣X���ta>��� ��op��gg�}R�S�J �*��W`PJ�20��+��������řҡ�CR������h��M�����ӧ����mfL�F�%���׿�l+�3�
�r��_ƏN0�ٻC3�hU���>�}��Bf��.uW_v���3�?n��0G��h6�Ga�o�x�6���0��	���>�w����Ի�o���������5�B�>��O�x����>s���gW43���cqSi�����]��� �,��f�Vx�g��He��*��-�,S�3Ёi�G9�͢i����3�����?�7��Y�W�}�VH���-n��+���<���TR��g&A�gV���5��5�xEV��<3�|4��۳{����_{����N�E��.U_�bo(�no=���h ���I�µ���8����\(5SW�� ���W�`���c:@-��id��Ȟyv��mK�^��[ʠ�r� �3�R��4�*]�e{�n��W]��|�V+���ܾs��p��nΤlֹ"%��[>�D�te3i������)~�rb�Ŋ�������|�>�s�4}p�#���z���<��s��m\���UB)W*��4	�H��<�Č����Pu�0�&y�;qpC�7	�����N����;���8���
U(� 	�"� )R�%��Ȓ���3���;s�{����>ݶ�n����H�{�P`����]� J�x�9�Yu_ޛ�o��÷�p�=s>:,����W�lY	}b�x|w��c3ܥ�t��`<���7O�a�?��H����5 ����U�\(Q'6%��rL�Y�:^�v�7N��SKВvs��ep��%���4K����O���ǻ��-t�y����Z����ψ��1����G���Z���ˈs������\��6�'�1��%@���|��K">����)%H��خ�86�)�FJߑ�3-��N*H&�F��zJ	ev�嶲�j�p�=�7)��"�����E�;`�A%��"��"n��޴�z�ߝ	�|T��~ ;��w��,���%	ᅛ�B���yj��|�k��U�9'������o�Xќ��߅����G��h�7�G����)��s�縼�Zx�0�\wj�؀MFz)�S�X�c$�]��ғ�e��7�}���v23�,��|F�sAV[�Uc�q�N"�	���������h<���e_Ǐ�[��8��f���5�i<Y����=
�j89m�ՠ�:>�1��h���fT+�����G�r���М�cE��1�`,�Ͱt�;���D���\���0����,Ǐ���6�~�����������n⸛��f��N�=<��bfk&3*��?i�����|�tn�v74��ќ�F&���J��̥�P��n�>��N�F=���~f*��\��]W�|�pQ���½��n&ϏJ���l��� 9���d��M�#EZ��U�՗>E�RĀw*��o,�x7�`���+�;~�T��y��R|��v��+�;]�O� ��d��]S'�f��ɝ
ix�l�4�C'����,��ah8�5��PN��ip	��!���[�Qz��η.�]K�g��ok�o|#'a�P��w��U���l��>y�tNU:���ɤ{x�e�V.��Β�.��{;��u���Oz~�f�r�`�}=hK�>�$'N��x''�]���o�ʑ�ǲ�}'�w+�,C$*��h:�p��d2�d��c{f2Sd?I˼:79����3�Wu�ĞL��>���钒;4G�i͋LV��ܝ����@:pN��ҹp�I.)�% ��1P�:���O-�ݹy�A��ow4����z��}�iw�����	D�T@L������^~����a�7�0t���4�i�x˰Ǭ��t;n���E��^N���{"���Ń���}�R3��Aє'�4�2��g���0�F��4�fW:1y�e<|���_���_?s��ɝi�U��n��������5\��SMaG8w��G��Ó��9�n�4�+L��3�y��I�҆nH#z���w5u(���B����>p�<M��HAV
>ib)_��V����Hw<�Z�Ν�a�/���[c�eQ��
KJF���9m�T ���t���0�<�N���x���SD�p��9Zpt�ſi�2nnn7�v����C����Ϡ�
[N��=&.�j���=���K�?}5/��,����������hcUSZr��x� Uٴ̭�-=�
�H���~jl�OGX�Hcu3K.��_%���J�Ѵ�whȽ��+��<���G^�ͭ�}<�l��(��1۠�S�Z�����4�]a#���V��Y�N�+��|�`~w�ۯ�}�0#Z�c꽟�4��ӈ�p�djy�=�1��x]{.<F���6�o6	-�Ȃ�4#W�&g��Lm=��D�g�}�NJ����Ȭ�n���6nϓ�}��s�/��ӹ�c35���粜�L:$g{�:�2���X��O�勿���vެF90�%�Jsf��w�d5�Ӑ+��h��?.ݳ�F?�T��1����~t�}��J���T��Y�pJ�.;�j7<y���84^<���;��,�Ϟ��/<�|N�z#G��Y���w�r����=q9�ty�����ek�&WL)z7���.|�\ґ�6�?[i�t%��B7m�dx��.��X��&����F���7���Դ�|�7�c,�q�?�(G]�Q�x
Jú0��hd]jJ/-�ݓvᇬ�!�D�hK/���2f�n7��s��\ś���gnw�X��[�ɖi�1�,y��97ݥ=��w�lxn�9�p�%�)0���0����4~���k�	]Yt�;|s؆�������=M5�2� ?[���Sh)�Z��z%z�A:%c@�xO�Vz��hDg��ݡ�����f�Wq	��ӽ!�į��L����:�·[�+,�~���0s��תc�0ms�w��Z�&2˶T��Nt:��yj\E�4k���b��$�r��z�����s���/%I%��~g��nӃ��R)���ۈ?D-s<�Ҝ����F�=ӊQ�Z��Vg��g�s���U��Y'����+�( d�(�z*R�[�&F�T�:Y!���P��A�x�,Y����ĝ����N��Z֦�e"��LkSfQ{)8|�_4�r^����!�Lp� �&���ȣ��M���M�a#��XF�-#�F*ƉCYޑ�]��c���w)J⌂.�q�F�x3�ԣ��
��)~F_�Wz��鸕#6�#$�K����s���q���F�����]˙���?
8��e*�ª��=px(�3y����ǀ�ȣ݇51�b�w�y��6ݐ�{A��޽t2�i��~6>��3�t?M�ը蝤�^�z�̭��<yn��SO/n�.���i�o�Гi�dI�b{q�ӛT��襗^�ݏ._��VmD�2� ײ$w4�9}*r�X�}���X�B�ys?�Ë�>��#��7o���jH�8ا��/䴠���>x�:/��#.�;�Ʋ.?']ι��v�і���܆��ߋ?=l��Iz:�{J�jȏ�%a*\�U�9�I��KC��$�	u�<�ul	��4����(�k�����ï�Q�kɏfs�텸?q�s�g�څ�ϟ?�x��'	(�8襬u?��K�K￿�����[��Ņ����2��~�����_�Y�k�\*���~�W��x=��徐����Qp�f����$Ǵ9qj��/-��'�c��ɽ!�\��,M��W��8��5�o�ҴHw�\�B؎.ٔy6�j^:���J63��@�a���4��i�j4o֨�O�x�f�^z�|���0��?���.>�Q��{.ne�v�Ai���K��CO�E���r�^���:i&{r�e��eS�4�H�Fr��tT>�w��J�E��t�l�7������ѭ��~�oR����A�{���.���8�����/"�Ojo��7���i��l�=}I}����l7r��G�_��:����I���~�1���t=n�%,�H��d6�� �a����+�g�1\\��廋}���s�2�ñ蜎�N�cɧf8v3�J'��L�,{�"Û��X܎���>�x��Wο�x碋%�L�3����͚��v�j��~�qw�;�,�2��6a{o*J%��dk�Vٟw3�R����yJ���S�A��V�ԃA4�n�S�0�r�A�A�3!>�i,�r��VO,yӷ�x�H�
3N�K�[�3;f���a̤&H}��?��aM�#���8܏#N��2t�[?5����x��mJ�pp�|���oR�p�&Q��ߣ�6��G�S�o�)��] �a�{4*����6Z�[��(��~�H�*q[�P�tS"srwF�~7�E�[k��S�<�߅�.�z���a{Y*H~N����C)O;�+�ۨ+��%DΉg�]m�-YU��[/_abF��`?�`�-=?4��7�i�Ԫp�7x��0iF�idm���袁��t�e���o3UT~P�w�����\���^q�<��<�?�{��$kn���ޛ��;��J��C�~:i��)��t��sP�5CQ0���(�q��	6���v?h�s��t&g�&L���HWe��#cz����f�h���|)�v2TN�诼�_�tU�5���̝��!#_k�`��ɨ:�4�K?旽)s=�P��༓H�]�a乂�qb?*������l��g+~̀J�Ö�����u��a���
^�B���S�ͪ����[�P�+udQ8�xq4�+����h��k��ŉ����qx�ßݦ�W���d����	6�Zrbt�4ܿ��/g�������i�����j_��R�B�G`��)8?�IMFY]0gY�������K{�D�}����?�ۮ��n��|�+Y3�x����W��m�Nz�q*��ޯ}��ο������e�����������_OGe4n�� V��y�e�x����`zkُ��h�0�u��xF�LWj�Cdw.#���֟��̞h<����;�Vc�N�������/��M�׫Q�W�9���l�2A˔��O�t��j���s�rq���s���T�OF����7�p�������K�W8����¼�}t��{K�,%���썴�4�)J����|5{9��u��F��򦟾y1}��JCG��_�fAN��dv�r.{���2%�Y���㕏��׾�q�y���4X����m�oNd��o��9��̓=
N�r��ɺtX9��o�ˏL��Ŗ�8��i��roD���qW���{���5,ljv��������/>��+���2kp?��'ΦCx��`��ښu&<ol�������$�v�4(�g;��n;Ry��.�{��j��R:�o��%Wߪej��}�_^|�eNwr�!��d�ͫٗ#�0]��$��m�Lx�`���Z6�~t��ܡ�F�����|:��3�'n��h~��_��^����O���c�0J�d�O�/D4�-IӞ�nDC����%S�UA�P����1�r;h���Q�9t�`�x����3��_ڳ5���w���r�iB!2���š�D~�k��77�r/={��#��ul�*�Z�+n�?��݅e~��;�y���%���K��4C`Zn4����i�O�[O�5/K����Ҵ�'���|�.�"���p�s��f��C�F��E��r�;9����p�?�i?6�	�0����O����C�w��l���U��FOrj��ܸ�s������[�5��w��ۉ���e�b�F�
�~m����F�AX�p0"�J�ὫP�����o�λ��� O�K:��ѓ��,Yo#�s�>�k4�~z��b4��"Hw?f
pi��`�z����5���k��`��gp�*�Ю7��Ы�"��}��x�w�A��h�������Y�t�ƹ��
ɔv��2�ˀk���g����\DC�ЇN�!7��Lx�0�b��fFJm�.~�=<&���w��sS��ڿa;l����LZ~i5�v��|��dI�׿o��~:��ַ���X�����k--�|���ŋ/=[�'�>]���?���6`k\����ש5:&Nv��� ո}3տ�˿�%5[�P{����S� ��H��ŷk��w��/�f4��fp#�.�|�F�th�����?-����U:J_�UT;�J^c�u���k���^�kx4|\�����P3G/>��34*���#jf�,�W2�O�����|9��%t6%���iX�sk��S�AYg�Ev�:���x#�nuguԲ�����L.#{��w�����b+�;�������'���or��nF���]��GYJ�5�7���y7�0i��e:6od3�����<�gDG��g�9��Έ�[��	^?�o%w� �l��z����۹���EzF�j���7�]�/*�._̐����>��]��2���-m��N��gߞί��h(�:!��2��*u,�M�h�������.�Ϳ���?s>Ǽ^�����x���U۽:HW?��x*���.侖�Q<��!_ȉg�S��Ό����s�e��t.u��������f���/�Z'7���y�A}5�ҍt�߯�^�����G��Q$3�R����i��ԩ�+�D8���3�,|f.��_���-�{6���W����pf%_y�eQ^|���-^������W�Q�������qJ&���� uK���i�ܰ�7��Q[-�%�r�p��F��u��#?v�����қ[�DUTl��Ua����Ѧu����]G���@]Օ0=d̔�+�D;����̇/�êNtF�Ӻ���D����ul�#Gˢf?�I�~��Ǯt��l�#2�,��_}�����q��t�h9�e/��H&���u�o�{J����G��yo^��M�w���[�����pf���<ޡ2C��.zS�:���n(K��%2�Qe]�>���_�2��'�O�A��������1�=�cB�͜�j�d�K�����v�.���=O�vk�G}W���L,K�U)�t/-�V��7����Q�s;8��^c��A��Q�X��N� ���S��p�*�	��0Ix���RnT_	S*?F���ȝ�SNgT.�(�%I�5��Z�-�YOG�PΡ�ܷ&:JNi��ǅA�4�UY��J��VU�2g��<��6�2.�P�[�~˂Θ�ä4�0#�i8�^/����A�?�X��6�jHi��O��ln�R�����Uf[�o*��Μ_0�<���>�m����?
І��iX��]\��=秿�J�(���w��WFW�g3K"�_#��_����{�\�a#��i�_��eKv�dN(z�翨Q�'r�=�֗kd����u�3y�d�֨5
n���,��_�ea���ۚ�cc�k_�|u:܍�qh��G?�[#�ٔv[�?84:�s���M�yА�r�{?=��at�uh[�,Q����~���1�I��8dД��@[:���wóF�F-�z�����,9�[�W���"k���7�����Af�[���o��eg���}fq����F�!G���+�l��[��oECػ�!�u����1��n^�e2�8�ә�$�t�EN҉pt�Q����*+zT�vFߥ7���~�N��IL:�N��N�N��v:��^a��e	\ܤ�~�@�tk�L8�i�5��b�R���1�cf���#�����T6T�O�8�&�R�i�k�3?y�u�98�����+��{��3��'�a�$ie�������3�<��f��Km-˒t�O���x�K>���(3�2[�W��ʷ�Ft*^���3��[��@Лo�|�?��b#KL��N�翐%[���x�������܇qc��ßG��L����Ǘ?IG���1v�,�8	Jָ}�Nm�~��W��������W��N�1�}�M��f�7Q鳞��S�'4��D����ԡ�6׈O�A�t�K�N���ͭM���`�p�������*ˍ?�tx�e��;v����y�ն�3�`|��A{��k�y_�kȢ��3��d72��/�	��۞��nm7ݶK�S'2��3�q;���M����YK��7S�6�E������D��o�t\В%�v����c�~a���>��ß�փ���>�����o�?p�p��jwU���4�.��F�>0��{���m:ޢ�q�������6��������k�ƽ��0�~�i�������hm�Ð5|���y�op�s������S7e�C���w5����?�����-C�X�8|�ܼ�x�JR�S���g,y"�����
�"��?��P���K����ʨ��#GiH�TX�x��g�B�z#k��s<����,�P�j,,�TհJ���P0�`@�2��HN\��G�F.��q�48hw��ϐ%ï�{��ʔc�v�p�6%�a���gc����0GT����6����oVK��5�
�LJ�N��ɫ��T�L+<7���g~TTp���������x:�A�ܚf�:�5jݔ-mu�<�c�W�W�Ͻ}�K�!p߄Ơ
������Œ(�P�k��5�pj�贘�0��M���5Xu(�`��{�>*�G���3��|\Yx���;��h�i��
���e2�U����t�pc�Ľev�6W�	�m�S������H�~��{Z_+Og}�8��u��n�B� �eD�g�-�'����~'i��	'�t��M���eS|���N�mg��M�n�&gF����nwN�Tڐ�G�u��d�d��a`�#N[f=�r)']
mi!�"Ղ��<V�<�)�k�22��Ѣ�Qn�=�t�{5k�cֺ�g�;�w����*#���y��^t#�@-qh�o�Gk7���I��w����~X�V:�Y&��H�u�t�ܭA�:�O��s�%��9>���Κ��y,=�ݽ����>��;����J	\�t��O���4��۶�Z��?'=>�-���0�`�?y�m}�w��N'u؟}N����P4�l{=铙�U.�7���ܚ~�rʾ_..�����	�����w�3kM�JΩ����z�˲0y�`B��iC?�4�vة���	�}r�+S��O�A���b�mSx�������7�0��1U��1�%|�-��TT��=�ݨ��Ƴ�}����x����o9����;L����>�}��a���M���P���d�qt&�mndP77y�OuR�!O{��\ʺ�3q����PuT�n>}��x�xG�ӱi�nÿ�������m���[y��^�G����s��N˫� |�ּ��?:3���9���Y���\�no�4-��q��ܿ�B���Q��A�y�c�<��!��m�[�!1�5�9��2�.`�i�x����sA���n��G*I�T�
d��Xn� ���:e4jI�"��Oh��M_FW�� �ʷ���*��T���1��Ր֘���(v�d$!��n�Ñ� n�S�͆��T׮�N����Cn��z߼W
o��u�.L5�m�7���-�Y����]�в7/(�� ���xa��C�0M�ƿe��B���wnNG1ꪁ�����4S�JFjF8�ʔ`L�O�-�|(Qn�<���'�|����?���>`��k���o�m��(�4K3t���/�Ґj�Ӑ��5՗.�ډq�l?�y讵�uI��Y��i?{{i��y�Y*)rv�x�T�GnN����^���w�]~A�y@�\���	�һ��چ�N���N5
���C��a4��]���^��Im9j�0�s���n7q���m�efXt���cW�v���u��������� ��4��r4��_�9N�B7��N�f-��M�0qN'�Ff�8��B:��NF4���C�>r�(?���v�����z:��̨4�F��-�t�t<u(ȅI�#߫J��Y)#�����/�������GA�����,��y��8�-͘�w�:����E�s�,��k6���n��Q8��+1����N�����9ǩe��%��'j��,໒;�[e�ƽ����e�[����IS�����şW������	y�1y��׵��6ep���l�:����:�⡃�q:"f���k~��/��AnO�K���J6f[w#��7�.�{��.�bv�w������r�:Ow�o�;֑(YG��^�;��V�2=+Q{����Ri$��,��H-���/��}��K�ĝa��]ǛzOX�6�+9fdɈ�t�U���6/5���O�
�6���{ �)�����	��3��ǟ�p�ZҰ�q��4�"���?v����3�O�t��M#U�1Ǒ�'�ȷ�TNi���W=Գ�gVs�y�\xcЗF��/��x�}�+K���H���e��4�%��'wn����5�ҁSٶZ�έ�A�8����p������3�l�1�iR���b��B���{w���O���3�; �ל>Y�a�C�����t0����78eU��sD�ixa�?
�p{4�)��2R�(��LU�! �m7�&�Z�U���eD�z���1àr4J�?u"d�B�S�x(��᪢J'������3�P�;�QW�٥�\�����9�(���^
]� I�K₣0��$5"35�u*�$?�އl�=��M�w��;-���p���3
���~�7Ӱ�m��;w͟���[�V�h�Tk�Jb?r ����Ę�Μ�ĐA���{�^|���ľ��p�v����O�uC�+��7�ܚ6�m��+~�S9"�n�k5��|���(��k��k׳6>x��gvH���IG��rt��É�CY��2��>R����D-��H��(�����8�NFߥ�T�k(��D��d�J��|��<����%��t�k�[�5����7��ˠk	!>,�`L��Ȟ[�����C�i0�gO�ƙ8i�����Y��󡡃B��:z�xٻ�9UK'^|kYb�g6ˊ��p�I1����x>v<rT��F?�G�G>9�+#��R{D�ܩ8m�(�jt��>��k�Bǒ�!���L�'�����؇�+g���,�����tCښ��w�����/�x���t-o�{oZ���O�ۍ�f��t��cS6�|LxO<����N����UWr9c�1�x<ri��'Y6e�A瘌���I����z���~Ň�p�ו�?���;�>����q;��8�Mwoٯ�r�H
%�R.+�=����	id!O�A�.}t���R�D��#a!���QN��IP�n_[|z��ґ.g�J�������+�'���aJ�^�d,/��=�z�^uX�Y#/V�S�,�J6�i��ܭ ��6��U�1�H���Jߓfd�Rp*�V��3����@]�GL$X� :�u�^�����Ef�8�L���az3��KO<a��o76#=4;����n�G��Fo��5VRl��-i6�8�
rd�pM���Vp�����C��<������2l�72����W����}�܊���8�Xw�$�����'�M�˸W���УpR�1�Y�z�D璜�P��U&g�xzBK?z��qA�E�GL�<����y�oK�7��3\�U���V!F��|�	L����x������>�I��w���t���;��5����i����.���If71ʭ���hF����g<��T#Q�y���n���i�Ńw	�����0\Ur�ԨA*��C:$kY�zc��Ѽ��4J���9�(��[� ���r�[♎�nF�2�J�jM����Tni�܎vټ�g#q�(��i'�8րB
GK<�.k���f�i�;�4w%�B"~*P��Y��9��.-��ၛ\ZA���Y6��XO�!U/e��YC���1%�o>��o�����De4���(���山� X���h�e��_2O���}L��p��v�<���;Ӱ��ڍ���kTf�F#�JȆsx�<Z'鹙K��96����a��苰h����[<��2�A�}3`ă��DF��z}�Aӽ�
�l�C�e���Z�<ɰeҸ�����w?i�����0����/��E���a�t8��t�'i7D�)��uN��N @��Dψ�����^��R���5K=*?h��F|�\�#���Mx�r��2�,�+�4P�!�0��tj��:C�É�Cp:���!��\����d��ړ���D9h��Ҭ_�	2z���(  @ IDAT��f����bu,n�Hg1���Z��EjK��nY��8u<�s��\~�u8t����&�{�-n����FH+L��pN(���k�^�S�`S�F�3�R�����
.6|�Kg^��Fd�~Y�������×��>y%:��ֶN��J���n.kY'��v��w:!��׮ݨ2�H��~fAb&�Ϊ2�ޤ�7w�)Y���xs� �%�LW�	�����$�{�bi��!�S~ihYnU���s	P{�؎��;]�b�.��흩�����[:��=�}w��}�C/�S>X����./�P� b:#F�+}��p����wn�]4�w2��o�W�����v���O��]&T^��p;���iHN:�|@�t��DX�Ď��G|������:��ѡ�<���gC�cn7_xl������;��lt<|����v!��w�}}�3cPn���Ж0��D�;<���Gǁ�x��c�t-�2jy�����ru���Μ��xi���?���U��Ri�_��2WϨc�,��Oz����:h�D���#C]$�sR��޻��w��O��g���ʙ"L�F~��{���K!#�F&�1��v�B��J6͡���q䞣��N"|�q���v:6�n�̙��2�F3��D!������B��̹�O^���'�;����Y���һz�Z֢���;wF'��,t�[�*(J3/4�y
v�z��(�?f�;\33{�X�7�~���dU�I���Me	^���o�FN����w8�����]�4�rZ:�
[#t�zp��d�-���j���[��FC:c�a�ҐIS0�;��vPp��S���/Nr]ʋ\S���$|��%��<���j�i4k���X5$}Ko��a,�4`�R�3�\#��T�ry|+�6����{A����,�f�iZFN��5��~��zQ���r2jS|例���*u�$���7�LK&��4t4ČzݙdZ����
l���	���]�����:]Qy�k9�m�a	H6A'��7��9�G|=���	�������T�%vʝ�	�%'���Μ�(�)�	o�/<y���H�m��NU�*��	N`q�=�;TB�����#��8_���2�%E�ދ�1`���h�g�����V�c����Df�޾���;��ws���eٌu�f T���Hzˏ���sXPNV|�o���^�hI{e�|�N	wxa<�,��R��W�x��F<��P�L�������HZ�D�Gd��/��<�yN������w�%��b-J���;�B���0p;� =C@�U�>�����2aM��ܑ����Ug;�V�׳�=�Vw�N�0UW�K�3��T���D�QZ�L��o�AFI�Ѡ������ї���9���YPU�.��t��f��\�:�w��{�>��2�w(��]u��&ѡ�G�/�c�xL�T����p0pz�q�L��~�G>����)T��;�?���R~i���^z76~��y��̲�
�K�I�8�p�?����	�Zj$_m栖{��;�źw_�e�Q����u������~��]zjp u"�hSw�N��}N�ﾣ��J�͓�{�|y�X˧�O�����g0�G6զ
B�7�������=V-��U�Uj�#{�n]υ�ٗ��䘊�$_aȫ:P�S�X����k�Y��O�-k����g��?��vP��,�����s�P�3mscʎL��<�)��n�O=*L�$ɷ���a�~���O,�<{&'�=�x��j�k���0I��q-~��;ٷ�n�L�����RI��GK�Kf��h %����h]$#~p0d~8a�T�8�7�H�9'f��Q�/��LN�{r��3O/������~Q�
�Υ+9��W�����)��b�t�+o)��E:�wyzRӕ��� �P�U�`�n��U`"`�a'�2N�:���([B%����q��V�Ke��Q"
����@�p�O�fm�Q��͵�״���w?X\|����Q�wKq�ed���v���J0S�7s:�����޸m�Qs'#X`���q$خ��|R�z'#����;��?=Z�ё!ۑ�����<�ý<-k~���G�|3l�L��o�.B���Ǣ�qxo\��Kw=uG-J3<t�W��BK�U�ѐk��mZ`ƒ���7��� ��w�����2�$3�"W��\�xVK*��ҳ��˸��6/�Y��&y5~v�8B.��8�Dx�mdtΓ���y�.Ѳ�� �̀�Gk��o�j	��[��O�r�O�߾+lx���|���aj����p:6���x����4�2����0�3*���6m�G�5FwW��W0│�w�ʟ_����ʎ;��ɭp�i�=s:�=L������ʟ���9?�yrV�ط�\pL-��Ȼ��wy�A����l�i�U�u�3������q�#�ݩ8���2�0Eczo��ȏ����s|������ �8��%�U�����:|�x}HV����v�7�ݍ���A^��t8�9�����k?�f�6.�����Ϳݼ�i\�=���yѻ��f�$�ѡ��ű�4��[x�4�����v�����g�C�T�iD��MN��]�7���8�_�ɔ{��s�����~��݆>�_�tf$�2���|�e`2~�3��?��R��e�W�I�*�+���y�MGc+�%t��>�`6H'Kދ���6�{տ�焁�\r�e��hX����k������^��t�/z�O��U�&�Е΋%����L���y$��)Y#���X�m�n���f�h;v��q����/�:�h���O���_8_��s�{2G�������܉��,�{����J����r ���[�Ymo]��sɠ�2e�/.�-��eX~��.��M�&�~̀i�{5�9�xxw,�+�_\|��_]�?�t�:����C����r��K�A�y/{�n��E�i�?a)4W��&�W��rFd�R �X���"0���b~n�U	>��N\9vl\�a*�C��bk�ҝ��۫^mF��V'�m-�~��:��hnɽ�����q��ȼk�*�xF�2�it�!tSq�3� ����:�/T�Y{&���=�)mʐR�7��E� �썴�+|��[!}+�K8�<x����{��cZ���~M�q�U��0�{on��tx���Q���3ב��d��8���O��i^�}-i���a��������k܍�X�)[s�r��~���s�h��1"8��Y/<�:\��7h�.�4nU�%�������6o(?���v�g�{@&�`�^�����X0C/�L�%�~��	7��|wZ��d֧�B#5)^<}�:��W��֨d�]%���H|�N-c� �e8�Y����ݹ��������P60�\�6)�v��Ѷ�M��!>�oԯe$L���_�����4^>`�t�����TT/݁�@�Z�ww�¤ȟ6�$K��~�_�C�<��Щ���;X�mpy�N"������۠�axύ���6���J��X	Od=p�ҹ��1Դ�.��gNw����1��m
Z��&0L?�R���5�<<]�^�0�<�?3�����ps�������"��1����+��,��{��=[4E�@��'�sN�{��7�[�-�҄ү�5
��
:0��p IN��|��]��đ�|�qoy��i�	QYs��ox8��=�C�M�^VB�B�l�w3g��w3˖EHGw���t��,�eQF�k�ԬB���&P֭��zu��*�]&����$gTc�LkrB��[��!������+�t�-��U}ϰ�����eI�W5�Un�=L��;��-��??��Mi��6�,�cZ���&nm�͍���i���+^-c���wVEA������Y|���~q�i{i�ݾusq3��yUN�$����Gӆ�>z,����C�o'}��҂<�yz���ik��؊[��L����K»2Q\�`�jVNI���t�.���x���\�����sg�kՂv�n���O�Z>�C%N��9������o^|+m&3fV �#�<I����m���+�f�忐�@"cdݷ5���J��H��KSDA&�Ь���p$�y
=�� 1�"����gXk҈���<n2=y�H�&�e�֧9��On,>��eR�f�v�h�"K?,[�/ܦ��cbS7
�2V�w�pFڷ"�$�݄יбݪP�}?B?9i��|POǣ�y�e࢓D�O��)@sx�L�U��o���c��k��4[J������5�~lޅ�F�O��L��>�Ԉ��P�^4��h�#\�~iL�i����@c�?
�;�`���q�{�ۇv���gU�����Fξ��Q|)�+��U��_�M�%ᆌW�����B��m���Q=p�b
��O�<�S��<޵�3��F�&h�ɤ�9��0�Ji*�}w;nWt�w<�=�W�k�:-��/������x�Nc��åC�g��R�u��O����9̞��O#��?R_���������(���O������_��h�&sa{]q�r���4�b�}b��3y��IU9�	��$��,�JG�2t�N��4g�c�����7thE�h�i�kض۽�&�7�6�<�f��#�v�aē�~�Y~������;����6}.�q��a���*|!���֦�ĵ���4�m��fn�έu�������2�w~���i^/�3�HtӠ#�2��c��'zS{p)O~m
>p+Y�d�|��ݨ����#ȇ���~�Cp��g��i�~��j<�~#x��� �Q��6��U~&J�b��#1���^e\6�ƳA��c?f��YΔ�Z��R�9Sb�w���##>�ʼE>��Z�0�v:չp�h�7|{v�z�r�8�۽��7�	���^/�F��"n�a���f�嗂�W����mF�U�?�SЃ~��i=���Y�z/k���ܳ�*��#���{*�ټ�����c��be�N�
�����A�����{9e}{k�ؑ'_L���gs�mXk�u�v�Oxй�����SIc�y��Ud9\��7�Q4���ܶZ�DI�<���t�՗��|~�'N/N�ø{�z�9���jS�]��{��'�H��Z%dV�1׻YJ�����������{y�)"E����8�ZI�{"��2��H�6F�Z��8��Jx��d5t2m������a�PY+��cǷ�s�)~����'c�&�n��P���%L��r�˨i�c?��W<���ϓ��I��vǓ��7>*��(�?�r1�,w�`����q��(�N�a�v����s���t�;�W%��p4o��Ћ��GwF��Q�FF�`�]w(:l7.[���g����t&:��cd�AK��̠5*����?n�����1���G����9=xe�����!����a�Uw~�ӽ���q�)�����޺���Z2ǅ�򂋑�ܛ�X�^^�⸗85�hiy�m�`���{�l�W~�N-��~������T:^��ͭh��W�K��?�NO6C�L�Q��?�o	�i�4���2m��L����i^���n��t�n�A�v��Z�_��̈4,5;\�3X��᛬��Ul����:~�w��g�,#L��a��S�I8�R���W�"��� �c0�������P(��h%1��eF���5她l�#�ކ��l��r�e <��ӝo�M��
7��_��poJ�|�jz�4��0샼����4����^�C��;����6nn�rc���� ��?��p�x�?�~�e�b��q�K�G�����[��0�1�H��ô|�Ts���6�os������6�-�h�������~�Ǥp�He�8�{k�gmG�H�-���n�xS�-A`�[;�����L\�?�*�r#zO�G'"y(��k�S�Jv�d�{D�*��W:)�Z��#���ApkP{����i�o�1��H�QNXNS�F�ɡ����u��l�����⾌�[mA�>",74m�h}ƟGz��倲�L�=�.���Lu��Ա��A�={v�̋�/�9�Y�OӱJ
ܝ�����hN�N�~ڊ	�8���Ǟ~*��6L:*�w�c�R���R�I��9}�����y�O�F���Ap(g�w*��l����O��4��,�:}<�I����7Ʋ��Z&��,)�� x�W�������o�]���-{x6� �G���0K=������j����n���HD�u����x�*�m ��z��<�������ԫ/H�pD���u�ՓO���	�/�KW��7�L�ًRZ�C�I���A�Y����Rh��p�I�R�4���Lz�Ӄm�^�˔���A���0x�?�N��Й/��� �;�`�
�;�4����?a���i\�x��p�Ԛ�p�U���*��~2'��ڻ#�� ��E��/2i\��\��ޏ�u�*,Jx��چ��ǻx)������[�̍���~�j/~�Vnߝ�+@:>Fq��np����8��)�n�jS��7�B�S)�7�÷���V`6]6��Ѱ��ل��gM_��!1�T�*%G��7��L�y�K8-X��CNL��� T.	�'�$��d4���t�ʛoޛ�m�IF�G���XG�N�=j�8���/y��Y�1��ۍ\Z6��A�x�7�@���l��X��q6O+�R�4��7����B�>)��R��*c�u:�hz�8��u ��;��3�d��,G�vl0`��vD0�
�|���	�ޤۨ4ظ�t���p��x��yg�C���v��<��9��)%��0#�(3�;���x�������n��_�l�����[��tZzW�Zv�X8<�
�+���/a�vw����� N�t�Q~:��2�vv��]]�~���w���t�c3��|�=L�����)��h7m��YM�p�Qvm������$�Q�#R8�#~�t�R�4.����4q�1;qV`4lS\d�!J2�K>]�K�����dw�v���m�c@��,�r��ۏ]�an��H:�럒�,4�g�����:5n*�е2e7���4�F�C��}r<y.%L#2�;���Q�]��VV��K���s�?���0 ���	~�Ec�zU��f��03���ۋO�\�Qڷ�рkYd@�)�I�mM��Hs�=�S'N.�}���t&�\�=9��^�������Q��n��|�}�g2����>��>X<�Έ�o��Ff>V�ܫ�x8-��^j�S�U�[qKi"P���Î��{R�R���ez@Ys�?D~�x@7�5��"��x����.M=afB����S�=Ws��n��\y� K�*iX�^�A�H�K�����S)<'㻌����B�UIU!��Y���-q�C1W
ՅR˯���
�K"_� ����T P�V$��h �{�I�k4���tX��#iY­3�������
���A�_`4<���fI��>�7�%���ް�zO!���;8+3Nq��g-���L��Z&x��+�7�L,�?w�;������(���
)�.��x�T�&��m�[���|�����6�q;���m4C��H����!�w-��F�r]��ϰ7�����h�Z5N�>�8�5�f�n��)���isk�>��^�8���ȧ�$��xz4H{��<N� l����� �zCY�N��+Et=�����7�s�(l9��C.�qD,Ӽkt�+���O�ei����g�ң��4��;��q�y�w�VF��C0Ž��#ƻ�[�K7��OG-uԵ#�u<l��f�us�J�lwL@�T���x'+]��Ew�<��iN�q�4>�~�Xe��ֱ��db�O:vxv匄Pb�?��/��W��|��e(m�mn���;ܰ�\-��n��5����7O?M���9�s?���m�e����҃��-��Q��9�[���n/��R��,�8�Sc�k�����]���5�b�|�Z �>z�B�A�0�%�ӽ�SQ2*�5*_��x�Y��	���[+��?3������)�޻~K�4�'�.������4J��M5�����xZ��-A��~zs�I.HU����%{s;u�vd���4˵�.�-eD����C�r��ѓQ��*m��3후͒i�^�Ճ=p�u"���ţx��d;d�'��)���Tؐ�o��{�7n�<#�
�a��9S���Z�8�[ז�a�xa;�B]�mv7Ky:}��)�7�s<��z�{���5���n�ц�[�����=J/<RY��\�ɱ���f�!��g��G�ީ}���l��X� Ύ��o�{W��೯E��ᑕ�ч�Խ���W?y/�w�=C�-ۇ{mgH��l�Υ�:'����l.{����c�J?���g�]��ǡ}\�|'�J�L�êS�(�<��p�	y߃m�:��yZPݯ�*,Vq3p�&��2}'2M�E_c4bNC�&e
=�-�"���o��u����U��C���f-/I��!��PB��d�41��`v?���'�fH�#K�ng�Mz��y���(�����;��
 3k��c|��byz���G��%��l|{�e��)�ݸ�צ#&��������ۦ;��2#��sd%��d=oP��T��g����~p07��uAMx��p`Z.(?��;Z����D.���Gp�Ǎ\���]�xաx�;���C��3�<tc_p���n4�C�)p1���m��M�w6W����������]�֩d�g�ס�~8z��-���
�7�P�)��7s߁x0%���.-����0u�B��;~f���V|[?jT�/�N��P���;7�V<�^��|ps7E��r����	�6�>��~�{�3@�꠱-�$k4<fH����s?f:Ƚ�/"����x�i���K	Qt�ix4�Sp�+]��ޕ3�'�w�b��$
��������T��nfN�쓤,8�����8�\�*�J����oF��6��ѠF�y.���̎;�ut+o囜r~�#Mt�y�?��5K�����0y��k���4l�n�C�A���3�t��#�7p��"#��3-��G��a|ύ0-���<������q�Ҫ�$�u�N�X,3���e��4z�B����;\�R�0-o�<^�b+���i�[V�_���,wO��k��w��p�6���.g���4�z��8q�ћw��?��rD˦bz�e�iol��sx{s���K�j�w�T4 �|*���GN��q{<ǘYL�����w��<�x<����q����ީF�����Q\�U��_�`��[ˣ��.-�D�<��_�UC&��o�9���BC�s�V��|��xo~�߲�ӗ�J#i1�!�U>H'���?z)�R3U{�����Q���ao?y$��5��(�{�h߸v}�ɻ�.>M�WmH#�6j�q���c*��s�'2 �B�[<��3�{x�԰;W?�x�<�|�a�׻�{����O�zgq-��Si.�gi��:�����c'�	���;wn_G��G�FYd�����83@w�b��~#�l�1`>7��(Q��Ϊ7}R�h��a�m�md�a�r	��L�)�|�t�� �9�|�~z�YǕ�"i6�(��+�ݍ_�,�fz�N��zN�z���Ց*��e�J���ز��B�-��l}�X���	�:u�۔����Д�*(	م)=���Vס�[�2:<��A�>��}Q��9'_��C�F+�F�XwI�>[i�)�ꢼ��`�y�1? х$��։ۊ*<w	.졌R܋l|�m;��u��F��iI|�f5�*	��x��k�L�)ޥk�P~i$�7@Mꔋ�ِ�K����F�}��A��[C�c{u���S��s'�f�I�.0�TZD��s�PG�kQ��/z
T~Ӂp���PJi/q׀�9�,�`�~#�i�O�?�FD�,e��5�Na� 3c⾞Ja=��1M���A�ӥ���15h�o��������N~[i��W8�G~#n�-�cQ)|qױv'���3��e��ލ�4�cw^������a�Vz,�%J��U�h=�y���{鷑��􎦛ř���K�(/�A��,^�%#k8�η��<]J'��c�#c�2xF�Q�����0�6KfI��+�S���?�Ocy��Q��w�M:4���i��onUŇ~<��4.��p�>��I/y
���p�[5�2R���9��d��S��jfc���������x�/pXrg�o�@G��Ks�XzPv����T��UE(�⭎�F�v|y4nw�Hs��� �'<?q�.���N�F���o���#|�a埰��?����Vd /z`��h�����t$پ�~�i#��.+�1���mԟ=b,�
����;�8v�Ttit��O�X��A�>>��A�7yK�|7�Z~d�1��;�yz͏��J��O�uƫpw�7��7��[����V�3�K��ïJV�5 _x��l�{֢�v�v��fy�^��[q;wSd���,��6��t�4o���)/��.N�����gO��hP�}���h�AgrO©�gS��L�Fܝ���c��cz*m����@�F���nN.���)��9M񃧑�J����`ɋj�I{ˉ�t)UZ�;`T�]�ʒ1�6s��x8��*�U���Q>$����!ۑF�2��+�F`��\����"�G������]\�x�t�����r�^�y�;��6*G���nګ�H�ԟv./6s�э`Gt��F6d���\K�2���)�_�lC�{bkq���B��7]��*M|�����#Y�t���'��^�ܾ��r�*��ՙ��ܹ�wo-�2x���ũ�ǒ���\~���4Ǐ�};�T��H���f���ū/�����s�)������6uGRc-�;��-͡.ʘ��:b��BS��T���TO�`5ު����ҳVm���M��@j�����r1	�.���$��D��P@s�Dn^�R7Na?�x�B�2�G�Ӹ�%��1��/��.�-�
�|�c�x�x�0��n�����뽶�,C6=az����'�
�4�Z��� Zʰ�JA�&��3�\�<���]!����KEr��*�ƥ�o�{t�F*�e�p�c� �܄�ʒ/�����[`�3��/��g�ղ���e:��ط�z�H�n���.���K�Ί��sO�.�D:�Fx�0CG������8���J�o�GOZv�Ǹ�v��n:�>��i@����������2�	'���.��]d�v�|`вy��5$���R'�Q��1�o�
l�5����~8/q5�N�
����Oq�V\�4m��h�A��G ��T|�����7>�Œf�;���l�C��A�W}��$O�[���!#]�3�ۭ'h����c��.������V� ���8�и��vġ�+^S�m�e��A�e1�`�/��ے�y�}��R�,��h������-��Me&y���D-�#?���0�����A>������d�����t�V:1pل	?8-��������i�O�gt�Q���S|�Qռ����O��r+��v/�B��Cx�ห7n7�=f��>w����)G�GCN��_#�͏�ǽT��1��^�Z.����\��Wó��,G��Qs�=��.��6�F�G>O��5���훷�&��L�����5�u,�d�t�ӊv�
�ݛ�_��oݪ4s
�K�]�9uh�����X�X-c�z�j
�Q�����I��Z*~�q�����!����r%)v�뿛o��q��Lv�~����)?����{n�����2�k9���by�"��H�ٶص�#b�H����K]��K��/�~����Z����`��έ�������	.����LN���N�{��1 m��>�>}|��"Ѫ�*72���c��(z�:[��NbԲ�>?����o~󏲺n�dr6��n�ؽ7��n�'���)�K�2��.��^�""��*S���a�~d�:��,J/a����M᧷�Ȩ*šD�q�R(���D���_`�L��h9/x��� �;�K��щ��A�#����fa-g/,E����Ow�v+c�O˧��ܚG8�|��]pFP�gF�ßI�O�>ɦM�㋿��L��!��5��Lǻ�G~���7鑰i\%&��j��5�h
k�λ��*��t�	���e	Pn�ړq�w������L˴�(nE/8��������sy���,�B��.�ܥ~=¶�0����o���a2��j.{� �Wu��kɚ���Ɣ>;;���~{;zyj�o� �*h3�_5�c������M�,'??��*�,�aLK��	��T!�A7���(��/)v�w,5ğ�B��$v��#w�p�\��[���f�,��![q+�r�ZNIcC����	M:ۧ�I��P.�4�'���}�i�O�����m9tz��NP��oy����Ȳ*���#`Z�G2B�v�Y�����|�����xF>jX��ظ;���ҵM����F�+�&/�A'�C�f�:-W<��GV�S����6�C���O�]z9iH��0O*�7�L�����jO���*��LK��y��:���@���q�P�8����7ՙp��ԕ1-��.��į����>d�H�tMY�,���x=�wo��e�iGN��2�ߊ�?O��_�r���c�c�-Es$_�;�v8+�L�T��m���ʩ9����^����O��U�:�u��YQ�>s|�X�菁��5���Ӡ�ں^�gYw��㎧������:��3�y?+2�}������,?���܎����g�f���4>�����,��Ig����'J�*��EN>���[����4���Hi��J��॑=^'7�VG6:w�D�y�t�χQfDK���Ҿ���n5��hx�FA��4�;�s��jO<��.&:{� ;h�@G:��"D<��l��g�S��9K�ϥCq&� �M���M�h	��ۉڃ��h����g,��E�,�Kqt�c�9��g���?�O�ی)핢׎y8DO^��P.�c�p%��"��6n��ą6
�r����[�7m5��F��C������������;�9o�$�����l�����sg��ǐà_�e��8�Gq�V����6�?>������ͷ8�a�2��_�E�K\s�����b�?���Op�-Z��z�^��ǒ7n����S�Pt�x�$}É�L�����9p���#�ӛ���4:��������eƽ��յ�Y�"�'���?x���.�L�ew<Z��FXO��O�N+���q?��M�Ӛ��� /Yțh�0�m8~���!Ԙ�	~�f�'�љ:��u\Іs�t���k�4Ͷ�����?w��1�&T�s�p�]a�n��?��f�4��s\��2����d�#��;]:���=A�]xp��$��{����'X2��]~b���%�r�7���8�&�aw�񁳖5Mr��B�O�g�5��F��� ��c�]���������^�ss��o�efr�ͯy�A��vK�7� T�ZN �4���{o�f+��'̝�Q��g�ͻ�u
�ғ8���.��v���o����pw��R���a�خ�tr�v93�ٍ|�~�ʑ��bħ���~���H9�2����
n�k˩e+.�a��:$�o�w�������FX�x븏8l����r��/~Q���ic�~���?��?�X���I�u/�H<�^�����r�]X�7'�|��P���?���|Jp������L'��+W���l�GG2Kqfq�d:yYn����,��n�Ŝ2��Vy��q��r�by����Ӿ�k���G�o��IK�*���Z>���p��{�׬��k��W^���3��Tڛ�;�U33�.i�f0hZ�Pt�2�!��p�lC�������&8��_���w"�ҧL�����w�ռ�o�a��J��o=�yb�d.�{,|�-J�Vh�[�f��4�c-��:4f����-Kh�+:�����?�OG�]O	 ���g)�Lb�҉�c��������"�yx�Յh��ܭO)x�-��)GL�㝻�5�}��.�}3`����y�4�O�%���L��0�?������t�Ñ�
'ܖ<���h%���+F���1��kH�OWH�l�zN��N��2�kF!~p��6�ަý�=�@[���w6�2����o<��8�4ݖ[}�I��õ�e�U2�l��v�4��A6jv�޹O�J����3x+�_E/e��������?�4�z�xx��|��k���o�'7n�M�J����3E$~��zh#���*l�*\h�CG�3��G�p&�~���*ra�������y�e7�6��A��s�q��1dr?�V&9X�h��d�k����xp�G�Ҵ\��{�?ps(�����ʠI��S�hz���[?ʿ��|tZ�7�;Oz���t���x�0^��x���!l �懗�aqD�}N5i��GW����_C�Q�1��h#5���厗�*W�Z��!��H(u�p�8��wǧ�Y0�q/��3��4�Uև��;4�\p�2W{�Pn~��A��_��<x<�	\�<|�BK�s
&���?��[C<nf��xJ'�ܻg@'+i2�k�B���#����Ox��|��}O��;��(|p�;�6�+͘N/a;������E�
���t�������+�Ӵ���h�i?3Kp��{m&���O�F�͸��f���C�"�P����M{5]ț������5�YZ��%S�\����鍔���8���.˚�3u�mzX�xcZV��i�~/�����l���NC��D�}4r�_,.mPz�;m:��˕��4,��ʨ���G����E�b$"�y�����!��,��B��y}Li�D_��L��V�|�$�ݤ�4�6�^<r,|qk��s�m .�o�@������dU�����4	J.H)�6"���0�M�R^N�`
�?�ie�o�-�O�-����Y��)�N?�8��㵮���V����<�� �32�2�'�
J�q1?qGCh/֭�s	tx3$�T~�?x6w2V�v!�~�n�/�2>	���f{��݅���h��V���v�=x�M��b��#�·�̈́�����>�Yv҈;\sYp�G�
�p��恫e?�m/�݀�T���8��Ž�&L�4Z
x��ev�.��M�y �y�o6����q�N���~��'����|�Co���ߣ^�7��k�Ï�Z����i����g8��پ��hw�[��5���0F��p
����趬Є���"c��(�k)ȸ��y��?�(��=�C������h&�q���t���`�����.Kr�L�2k_�z�Nq$J#�X������/�#kF����z��*��2��^�s3*�䱎H�B&.��c	 �@���`�NaÃG��0�Y�.7����nih�����4��	��_4�<i�trU�����c���ml�̭�h(��WnH�De�G�O^�e��Wy�cPy�#�<xo��#w���������S]�Wf!8n�Ӟ��]��sxБ<����i)���y�f�h'��F����Ǽ�:�ʇ�d����r�+^�OWۮ���t�!�'�)��Jν��[V�c���U�������ZY�c)����o}7��3HE3@�F�K)�liD�f�(��w���
�+����}@�	�_� �^a�ŋ�e��9��&#�6�h}�G:�&�٢i4JN=X�L����Zq����~m{:�`�m]�k4�E׶ҭ�E-em|�=������\��l����{��':����/���˯��d������mSw�G����u=�6��k�ڠ�(����¦�a�{�G����k7�Y �neT�\�O��s���i`�o�·|3��䋴=�r�d�=1��:}��tJ����4u@�qv�$C7���X�N��P��N��%a�,!�NVDGz�'�;�� @�q�	B��5��v���LR�W��H��[$WW��8/揣�h�wck��P�Y�k�V2H��>���H;����b$/|�Z<�;��<i�^6�������N�-J��  @ IDAT�����['����4(������!
�H'�<=ɠK�]*��H��4��N����� K%��T�^����(� #sC|�+C0�g�e�$]�c�K۶��sU���W��+<�"�4��L�t�T��-���k��&��g?�Vz�W���as���7��I�I:����A�~I�N�$Ly#�&�����<y�K�[�q�1�FF��암_�N��u���m_��,N�������K���H�6���v��p��_ۏ�[#�v{D�5�檣�|��a{!�KϥS�LGY:I��v��a[�_���ҋ�ʟ^�3 ���\w�3zm��3���]n2��Ɂ'Sz?��: #�|�^蠅6'~�K���ߛ�~��用�۲�r^����f�(I�����O%�}�{i��d��]���JW���?��#Wa����0�P7�:m��b�&�G����#0������}����]E��`-�=1�ۓ�g�̡��?���ꃺ"���u�{��ތ�Ӣ���R�1^�h,��;�z�	EuB��u �s�Gx��IkY���N�E�8��=׵}�܃�+�k� G$f;�S~�xi�P��g�d����m�S�W:ޞ��yֹ��w#������K��HS}��_�M[��g�¥߻�`t�o6e��;ߴ��ޟ	�k��v��C�2*O+��+�H'o�rei(�mK�F��SO�JO�:�n��Sxdq�`'��G'YGO�������:W!W;���M���^gy�4�ߣC��C.y�[&�y��OO�&)��aєs��y�V�L��p+}�Iȴ�i*����>�U��;����vrdR�����~3г�ԅWvRRձ!��w�ߍ<����[� �I���!�2�z�6�Mڎ��.�>J��_�Bɭ~̤"�һ7/�;�LZ虤��y���ϙ��}l#�Un�^�H������K�^�7�V]����G���LxL*�t�w-���w�Z���V�����E�� ���\�3�	��0��S2vx��a��&�@�|c�����^�P��l'��k⠯��7��u~�,3��N�d�q������y�U�)��_����GG|uL�&M��ӱxW�7�&�hֶK�U�+��p�j!x!t�wd�#0�z�k{�	w���_�V/��)��;�S�[;�<�Ŗ�x�K�cx4�o�_v��B�k���hɫ��$�l%J�t����t��P�_�-�<��J�.p������;�ov�����1��6m�V�+?���@�����h���1�:������ N�AÝmurdHc`o��S�ʓ�K��\���^>����e�q=Z�����Ũ�~W�Y�nu�zT.�.��r7��bF�Y�h��cBd�M��3��.�y�N+�zX{�7 ޻�E�����Ė��Nnvz�
9�t@G�My�c�#���5��������P���:�W�/=�������/߱�v�ǫgB0ډۉ�.����[y��*�]���W��K&��E�#�pĪ�}s���`k�^�)����KO���l�廆�&��LG�]^�ؖ�o/u�|�\���n����*�Mip��n����-������Eqe&_y��{��w�~�}��F�$Y��E�'��L�3����`�do@_�����Um���dB=�߁G0N|����%XN:����/��x�N&`K�=]��/]?�qt�i�i���\t[_�_��kk���z���;�S��5����YA�.��­?�}�9�.}�|��8agl���A��	Zr�.n8t$����ۇ�<]���f�Ǩ_�s!�;<;ԎQa�x�d��E��ӌ6�� &О��9�/�6'݀���W�w���� ��~?ۆrg3�z�x���2�ޓ��X�������W��S��������-����X�
;%|m;#�I>]
Pb���O;�y�7άr�s��Lz�i����Ϙ��O�0���>)\��,��a��E�A��4.�82[����<��I����)�Ӭ�c&�r?�g��X���M���N�c�o�L!n 5��ĵb�AZ�J���X%��}ȋF�#�QT$�
���tR��r���<��_���M���Q�����?� �i��sDe\> b�>�N�_�$���\|�U�"�t`�5�v��巁����_�~q��n�]�pw*�t&Vo� 3u�O�g6w+�Ž\�==���2�U�U�x��##7�D|��|�TV}��N�i*x���:���9����3�/��u���vy߁]nD�qV�b_0ݐf%O�*�:�8����<5�<�s�����i@^���:�܈�K�X<ۓ��$r�/8��Y�Z���$��4�yY:6��	�v-o?7?v��
&�d4v|�΂�����|l����t��;M~���<GK��K�/l'd�D�j}n+Y�[e4�Ь8�F�Q~�����&�_t��3��K쎶��>��!v�ݑ�&�䰹�)�̴�
_�h
_�����N��I�r<� ���Q���X4��e�۲��j�/��V�l�]��l�|�N��Y@w6 �����51�C�Y%�>���F��+�[��А�S��}�V�I����E��I�Z~�/+�-'2� ��#��%��1��F��9tG��-����Wgk���Å�m��r���T��AC�O�v���|�Q�#��z�n���O���eG4�8����O��Q��|Q5�M.ݖL^ U�����nĥ��X�?��#�������u9��2ue���a�SGB_=b�4�(6-q�V&�r�5�h����>���elF��?O�����;�m�oc�c �6<g�k�Ѝӿՙ�m�j+OH��t'�|��om}��3gܧ>��Ӯ�DӁYB�,�g��{���>�/[a�7�^`�[�v���������/2��>T�{��_�i�q��ì..29j��>)t�mqD?����n���l��W_�6�ݓع�P��K�����y�c(k[��s�^�O�U٤|
���j��mm,���c��S�.�1�i�"l����C-O��l�݋�V�����,�*�r�~��M�ئ���K}�gq�
ڮ�.�Ӵ |�;�餬b?i,���R/�%�Ov_�y'[�J?����0P�orb߼ĝ���;�p��'���c�lz�&c���� Y��{���W6�I�T7MǄ�իu���1c��Q���.��C	�8v�}���g:li�B �>�Ξ���R��)�7s�pt�7$.�^n8��x�n�D&�CӤ�$e�~�I;���oW;� �޸N�LCI��xt�ρUGӰ��x�	����O8���,��0������)�Sg��A�8!���rC8P8�A:���<U��b�F�I̸0��0��Y�[��|��}Ɛ����oZlO(����T�߆C�7QD��q�]+��1���?���y�S�k����٣�/~�$���A���t5�����x��: ����kG��!��fY|8����ÁǁoG�?4�400���3��//�K���o$?��M��i`����v����6[��d2 Ց�'�pU�%;=Э�d��<eh���D�7�Lc�X�3��\���k�F�-��|`�GOH?e[��<!��I	�n�S�x���|2�/d��*dB�<�ki�ꭈ8�R�<��*7�e@@v��¶hUp��C�|*K˿�MF�����|~��vݒq�S��ePa���t�|i}� ��Og'��a�ëCc�L4\O=O��V�ٌyr�hovC�u~&T��:�[Y�������zZ�\�Y+:O��\�Qw��o�#c�6��]��<�>�K�������Qv˭��G� [������ǐ\�����s�o[�i�3��M7<���K��x����L��F6�[]NM��蹡qpy�^m����a��Fޡ��+����T�З6�ɀ�ӟ6m�%����n2�������w�0��&����)��`�+�NZ	p��q�7x��7���M ��_xh�ؕ�p��zt՞���+�'y�t݇���K�^���Y�>��3Π̖E·�ʻ}<�p�P�����s���������;M�z0�c`o���u��_]��(��E����I#�#{7Y�!���6�%'Xx{��ȪE��֖��EA��:W��a�\���0�L�2y9;�B)[d1�,�K�}����0��sR���������D�j�ҕ~�~�=ؽ}�0����`�����/e��[�ِ��Ӊ�֙�����zk������bs���,����}LL��Y$��w��r�3��&:_yi���ɉ�Df�AM����%����7������������"�[���6un�ӏԨ��39�i\l7|���Z�)=�Ll��?��$c&��ia@�m9�*2]3A�#׉�t:f}
"��������Փ�_~�$G�}�	�7��f���/���Z�oN�c�ُF��o՘/����C���n�c�r�%N�oG�4����i���A�t��40���
U�Y�5�����>��%mu|kW�⟊�$�Т�\�������4q��r3ӝ#ł��v����B�J�\4iV�����C�kU��ҝ����j���N�%W;0ӱ$�60����o�n��	=�|\��ɱ�$WU&�-�N�Jo�v�,��Mn��՛
���1��Õ��7��W]���o�zs���_������2��Z���Pe�H9����~�&����U𫞭:!=DF��Ox�w:�M��^��Ƌ�Հ^u�=:A��K�d���J�z�v#�քA�Ќ|�qF�~����>�ޑo'6[�����AXt�:�f�� ��S&���co�#���u��*C����T6:��� S�)��o�eh�N0�����=O4Zg���L��i�}W}W���g�9�o}i�px�%����Υ���Z_�3�#{���0�Dc�꛰�BwH�NGJt����/}�}���]d;�<���I��X�~��������]흮���7���Tۮ�M�=őϑe�m�Ypկr��gx�_n�2Un>�6^���A�knd��x�g��4�7i){<ຆ�P~��?�L �<N����l<u�<��%mmW]����$�If���&\y����k���gO,����6���I:h���]�ab���z�/��-�u-o���{������L$2�����<}~�ck���W��_���|������t��~��e�їkK2�M�]��y��-��V��'}���~'�5[�|�n��y>]����H����ɣ{g�9�0f��ΔO�gq-v�4��Ө���>OS#Bo�/}B.���h�X�3Yĩ��|�M������U�د'	9�)�eD0�I'#��#��o�����Lld��c5m�\��%�9N(�7�u��o���4Hn�S�~˝
���d$��<_dU�]�~��p��o_|��m{�B���}C�u��n�����8��h��-!�z̹��or&]���9N'�у�ve£t�q*4��⤋��o*P@������}�<:�m(�Q:���FVp�^��p7yͨ��$'�<��8����3��$�����\et�Je$w:a��Y� ���e˂~���f����'O��2�VV9nd���4<��<G����^.p��� ��˖��rl&�ȭ����L���{�)�y���`�Uv�����$�[\m����)q���F�m��2�Y�^�\Z�g�?=��?>U��ܔU���'e�U.����	w�om_�4{�����/����{�Zr�Wt��o�ū���*[�]�TZһ�a�w�����.���x�� p�Y��z�/L�\��o<^IZ�]�/~����:Tل�_�V�(��N(���kNڲ�*_��O��5�x��v~U֋F������Yکzx�=���*.V�=%md��/��&�>|G��w7�Ce��UQ'�iٗ��<��H;������?r��~�Gz�<�.^��^��b�� M����`�k��w]Ͼ=	ݑ?�M�lt�E÷���18w�~Vz�N4�#����Z�{�I��y�|��޽Lz�;��-�����A���N^���O[�Ȅ�l����e�F������ q*��ז���UΥ���[mC:Gz�#����L�R�Ϟ�d2�|�y��O2�x�oQ��9?|��|��;�;����{�1R���*la+?a˗x��-LeJd�ǈ�o���_��%_yVG0t[�~�r�.M��?e�md�y���YTۗ�׾��]���#������k�`���}���2����H%��fvU���eB�����K��d�GM[/�o�me�}�=x�y�T�z�
�ѭ���IT�]����f$i�n�dք�R{W~�\&�"�^���7&������9����N�*�������S��̄⛧O��2{�G�A��b��i�ٌ+m�1���woA���/y:��u����αb&AY1B��mS�*��"�p��G{=�:�4~_xD�9���yfOwh��䞲�祯�	�Mg�7��0e.2�MC�=F��V��c_�ȭlG���%+e�zL��l�ʍ�t��+���M|�e��uS��<��_��˗�À��<���58�u���['[=G����4�����#��xy�EN.�<ݣ��o��a�	)Zl�6{`��I�'.�u#h��p�KO���Ȕ��}��u�\��30�����r*��Gz�M����ea�)��tLG]j��Ǔˏ<}7��v�Z庑�?tK/����ʻ�W�E���	NG�|�u�
��!y��p�.^�~hՅ��	�e;r�>E~�%W�.3�_u,<=ѩ\ss�T��w�}ni�\eM�H�cyE�� �|��.����e�����i[x��<����>���7��AV�����B߱�2��l�Z�P\�|̉��0#)4n������w,G��S�Oж�(�;�WM��@2�7�ۙ@�92�UGj��bx�&��=/0g9�A\��/3�� \�h����GF�o\�������[���$��G���}�7ۖ��=��|���P��.�A��,`�/m/�kt��ù��ŕ.����:�ӓ��V^}�Щ\�0�����h۰	
?��l��Gc+4���`�ʋ�j�M��*��vv��������E���>�~�1��r)�;y����Zd;�K����=��ѣO����~���O�e�loM�$+��mě�������6 ��}������W���Z�r��³C}�d�16Iy�gBy�1�<͈�f1˸-m;�cB/�w�����������9���������Y�e1c��Xp2��D��H8r����g17����B���)������I��(ntI�] i�I�m��s[���z7���r�KK}AS�0�󢺧!��	�JR7q��+m�h(mj}@�|r;��,^t��4L'�&������EЯ�~~x�'Orb�`��S ����!���!UH��ytK[~i����ȮS�)�T8��<q��<��c�Y����1��ud�.e�P�}�Š�����k�Hejz�H�][���Z����J�*<�&-�k/0���0���X��^csn���b:��N̙��a�@9��#��m/�8W����l��eW�C���~Ȥ�٤L�M��妁p����Gg�+��V[��6��� ,��}�Ҩ#7/�_������ћJ�ʧz�?�J�q!F^��.�t��<G��4�0t���h亸X7+y��^>���ʅօ2��CW>��	�yhZ��Zü0Y�Qk���󸕳�n��t��[�{��}�I�UNaȏ�t��<��.����._��oݰc��!�/�ĕ���:�љns+�*g����\�u�5��ŧ:Xa�.���O(�q�
㺼�מ�Cj��q`���,����'pOr��<|��]绞�Y|Y67w��N�>NL������c}_R'���|�]��L������C����]>���枵l��z���CHN����&3��M>jF\xc�b�8��_��t�����/�+��hˎTE�,#�6��T%�OZyͻo÷/a��Z�9���K�����_��--txy�&/R���ױ��I����@N�`\��2�g{2�h�.b?8��[�M���G>�������`��W������zyd ����D|&�Y��v�B��w2���G��ٲs�����ɳ]�¦�Y�˻�k�����ewu�����,ʁ��r��nʌ�:{ٱ�L8x)�y�$㐋lq�p�	��I�mʡ},~�9f\�HM���d䈭y*�v�7�y�r�>ɋ�7n%'����\d���)��7�~;`,~�rop^�)�]܅��xjEDZ��o�o�����-M����XS�'2���.�7� ������Z�9a����7��p���a5�IDn	G94*y`΢�'//N���ċ<�ph<�W�sZE<�p��6E�Y3�D�`H�5��0H�o`���Z�sJ��m�������}t�p*��UX�L�\*��lelC��s`w֩:
��Ȗt���Ɩ[yV�����qH�.ل�@�=�寣����ȱ���]�]���4�i���� ��K{^r�+�͢�J���[WLH��c���#���]�Fgr��MEG�0�i!܏Ei��N�_����M�֦����~�Mi�囎\�E&�a�<�������X+ZKG8����Sm�W��0\a������׎`m2Q�t~h��)��uVgk<�LY�=+i���>����ϗ�2��Y7�I�<p�E���S�l-_��8`���^/��"gh�̧��b��2tW{0p�C���,Ѯ�O�$��ЯN�ށ�]���//o�M�ܺ>�%2��E����}�<�ϵ�������8�Ȑ�yZ6�X��!N|�C���S>`=u���iCl����Qv�ya�d�8r��oR[y�l���h����l\�ϒ��DHm�7!և�u��I
ݴ5�w�(T�W�_�h�s�A�t|�Ҹ���#�o���/|�y��������C���:o~[yW�n�ڠa��b�������9A.�c�?��Ƀ������]_�����|0��W�uW�Fqy�Is��Od����t��6�����+]= �/n��+�@|l�A����]���?u�刾�o�W<!w�Jǧ:��Kِ	�'k^�=I���4�7��>�S���������Oϼ�o���i���D���p��>Mq�r��v]���oɸt�0��*o��i����S@�x��i���"�ϼ#��T���[�ɇc�U�S��W���F5z�����Q>ʄ|S�S�s��8�C_o<*N7A�ŦL���Km���0L����j��^��44�Y��^��XL�^}x��)��}�涖�uq����w�C���tS�������[A��S�6jf{��m2�N�M|�)<FS8�8��Q:ҧ �_�%ڠ�6l><{4�=2Uat$]90`����@XZpt�u��"��ѡ�z*w��pOȦ�Rط�
���p
�n�d(24.4�w\㼋��9�v֎�-�xp#Kxp���V2�i($���4;^d�Y9;xu���Rr��Zٳw;|q��d����p#�#r�VFx��K�t�&w�����H��4Z:�A��^ܚ��N ��Z��9���k#�{��M��o�঳@�,����ny�c�P>�z�+Z��Ǒ���֟����
����!wuzpѓ�n�֍l�K�Y�� /7��l>w2�AwV�"3xn�`Z���+;|n]�t��������-j8���'�U$����{Z�	�����^���86l9�F#Zv[t���Xz�v^~�Gs�;�ë<\w������ƾV��Y[/�Os�l���[fhù�=e�٤�ꂕ��q;����!�K�U��$�s��Fc����-�zY��z��z�YE��l��K���M�������7���5��[�߼YO`���Mf�y���S�h���B����b���^#Oh�m��_�V�6��9]��c�=�s�o�����"ܟ����w�Z�"/��ԙ�h𓶵_eN^�y��5_�����ȧ�Y�-;��2��>�����db�	z�|�����7�_>s:ҚP�KN�|�w޽pd�*�t����K-�G��r^e��r��4��ʫk��v3��Oiɧ7>�P��O]�!�י�}������ã�/�������g^O��h�]\�jCK|x��u���,^.�%�����%#��$�kz���2��#N����wߴ8f��84�31� z������I[��+P>���R�S�W�#��pw�`8'%�.�G�L4�Ӯo���7O��L|е�"����'#O�M#�qܐ6M&�-�u
t����/��U��>@�wy?�X��ǟ}���Vڜ-�3�1�ك�fVG�P_��ܸ"�i���Ǐ�������'��r�O�M�ؗv;�a3�� �7��e9��e��ّ�'9{�o�07.���Վ4��L��b��i΄G��ƛyD{7��A�j(�p��L\au����裏&� �t|;����2���Ttx*�*t�ޫ��&?��ro�h����P���W7_gH���o�龏��t�T�`��\a1�3#��@y�B��O
��:J�'is�^m<�nK~�*��+�2���ܭyg��RV�R�C+�We��|H7g����A��ԗ��SF��������^<�䯍�L�[��N�ّ��B�9�:�~�{�&�s�l:�9�\�s�n޻H}v}��A�6cS��2�lV��ݺyo�\�Gx���_*�_I|���5ftqx�Q:��Z��"���;�]����ҕ�k��Qڵ�L
��T`�D��6�N�F�K�躞�-F��W�����ӱ��X}<�|���J:�y�ܱm���%[:M/�Gn��u3G���@Q�"�mx�X	��0�x���U�ֵtpB������~�'4f�f���FctM��*^�#�z7|���h��ޥ��b[s�8\y�r�,9�'�C�z�����$��}<�0��e�ͦ�3�ңui�3�M�p�h_������(0<�zt>��3 \p��%�79��~�S����I>��l�c�w��~����o�:|r�G'����ߺI��=$ߤi=�;���+<ғ�_���h��-/�V=��=u��L1v�حv�G>�p������}�>}S�S W��w�N�}�9���q�>��L�S	R�Yز��>�U^����f@�24���Xqj�<�N��_�u�	߽%�,��&-�,���G�����K��^��~��A�ׇ���K���-)�����i��N`_�|^��k�Nڙw������zQ>���{�{������\�0q���ō�+}��ʮm�U��9�@>�oZݏ8Ug.������# j�oS��Ǐ�3���_=�Z��,��������1�6�[m[~Č���$y�1�[վ�� �gQ2��,�8�Ɠo_�_|����~�eޛ�}�⋜���u���y�S��cr�q�B��k@I�i_��^\�&~{��C�2���}�?�s��dXm:v�`��mS3�p�٫�o&�)p}�XA�I^v�xړʜ:߽�/z���1�����R('{Γ���U\)Ә�,�k@'g,ʽ��SꟅ�T�Y�L����J�f�9}�����0�`�}_g0�2���΋��"��#�u�&&~�^&�F��l�"����4㬜9��e<��E&�Y|�{kM�o�~�/��|3q6 ?=�"q{��g{��翈̷?����_������wmO^���"�oPX ]w�a���*��~WS �E�T^���3����W��9�{���pAK#�n :^���q��&�����;��GS'��o:�\�7�C䔇z��m���z��N*�38>hr�G��)�h����i���-O�A!Hp����4�2�|i�F̓>�7Y\W>�8�-�҆����3�4"/I��{,o�\X�I[7�e�$m,�2����W��P��E#�p�:���C����|nN�1�5�z�6nd�m@:OG�TƑ'��V��X�&wp]�}��S��2�����]�S��K��ʤ��Z��_��|t0#��iMՁ}&=
r����{�M��i����k8e=S|�Ϯ���m�����]��y��(yu�at�u{�Js�^^���\s�Z�`٧�rd�(�#�:�{���ep]9R����6!D�n�\�C8d+�⻾�O�k���V�n )�u��S�����+ou���t�<�2A�F��Xg�R]��Щ�,���t�t��C��]����Pw����+.��P��ohՁ!K�K�������8��p����_Տ$+|�ߗH[}d�+G��d��k�d�����S�]�K��؇���G�U�^��$G�Vwۙ8�&j���o�#��֡�9�#"����'?�?�����i���}���8���~Tt`[�|�'����<z8�/�.���wzj?ai8��|�q��V�n�"�ˤ��L�V=#_<4�~�w�3�d��N
��2f�;�����~�q����q��͂��|œ������� ovp�g��j0�gMz��L�h��6f��{����I ٔc"Y�L������{]�Rf_��Ë�i])���U����bN�neb�B��!M~�N`��ݦ�j��.�o�+�L��u/O�,6���m�gd������u�����?;<}����ԧ��`}����o=�!���裚G-��wݡ\+��6[��ud�`׀���S�1R�9�v/�Ѧ
�MeJz;0c*�v*��[�V'�,d���.y4��#�:���ި�QF��l�;�d�C�+��5��@O��Iņ'^'��7�^�
�po#i��^Ze�΅kz�ˣ�G�d�Ӫ���P�In�I�?Ocz�_�1.X�
������&!�n���>��	O��4b{0�W���Oy�guo�qF�ͬ�<
n�X�y��lQy�˷�Ūk�f�[R�&���^�'/�dFOρiH�*��ڒ>d�Gnt��U���ө��{jY�@m�sx��8�Q�%?}�Fڔ�'6k A��S�	���s�a+��{���c�8y�Ł����J�q��M+Neh�k��O4.a~W;\��I���n��bn\p��r
�'M��:��]vO'��:\a��4������Z8G{冤,��k.��6��h�<�|���b�<��Mß/oq�����ꏴ£�|˧r	��]��Z씓��f�ޔ}
��o�Ccɼ���Լv<���o�r�,�'���M���M@���h��^Ҫ�tqm�����>�hT�k�l���-���~|?d��@�<�w�%���p��șvP9*���zW7�k��ǲbs����� �.`_������{�}������v�oK�Ew}9�}�~��,YW�����������8o"j{ѽ��W��*)+�,�d�)o�G~:��	Cd�v'+ַ3�m)M�^��꫆��C���~r�ۿ����ߌ-}�����C��g/��+O7�?������H���vR�c��v"|��g��|��ß�������v�sV��b���~v����	���R.�E�V��ע�e���Y�m��2�I�re����z�|�Ԍ�u���9�.������8��o���8������O2��d��N��%4���2�����{J��4�ԙL����������F����6�ގ�2��=��� �aڪ�w��~��ǙD<8�}���$�*?�������蕇r[�]��S���>]+�4�X�5��̣�[�0��5~O�\ĭ�
��vp�T
�G�u���A��,*�T�-}�i�a�Ӫ��jh���욬<W}+�Z�BD���n)*|i�eG_y����8�@�̐����G���M�^��.�?x�7![��i{]���;6��+O��O�q�w�ڄ�<ey���N�M���ц<vO��>xh���<�Z���'���l7�p����g�����6���I�
G���G���HkK[�W2V��ȯMK�y��l]m Ƅ�|]�[}mS8ʹ��.�W9:�8��o�#�/�+ݞP����l�a�>�>ʬ���X��Uw�]��{��-�"�eX۸��)-idܻ�%��'>��8��Pza���_\:��&y�JO��ɍ��K㘷!�]�-<i��qE�27����-2�ᥕ�\������5��?����/N�*�t�L���a�ʨ����E�s�-�WM��ϼ��:j����ܛҜn(�N+s���m�i�:���������U���k��rpx�����F�����n�����|g��\ブ�#wEw��/�����o �`c���Zf=ݕW�/���-x�Y_�^}�w"F�� 7��xq~��(��+�U��}��@uF�q����@}ig��x�%5m�����eyd����t����y��Hx���Iбznla��-wQ&�����%g���l){��Y�/ϟ~�<�S���n��#μd|��M�l�x���B2��|�yc��l���?���p����:���?=����E�(�f��	���������H��`�=|�Q���b���is�L R�y���A��C�xm睢�K[�<�H]�fN����{	O2}�3�L���>Jٟ�����p��4-��,}�lg�'gbcK��7ϣ�Ɍ'n��|hy�'m!x7���Su���ׯ�W�؜FvPx��ּ��"zrx�Qޛ��;�B����8�Jx�v����?�k r����
�3�oGfo�M{�4�a�b��vBQ���!qB��W'(�u��#�4���])hg[}���y|,���#Ge�N.�SaJ�0W2.������(��A<��8�"k���G'�h{�d�n"s�J8�P��{>�ǯ��Mǻ��	l�����&�#��ih�;Q`�B`���-t��d�Qs�ѷv���qe���v˻!Zx�MXx<�1�m�c��j�:� ����x��/<����l\{�m������-������-�,NMܓF_��8چ��]o��B����p/_y�Re��瘟k�m���g�W��6�r�}����Kz���ejz�z��F�n�ߥ�I�F�*�A��~��,z�J#k�X�&�˿����uC�k4�0hH������n�p�����=�w��^uqm[�4�N]ހwx�~�����Zq��� Ǟ6Z\�V��5�aen�H���Y��'�*|Ok2�"�J����^��[V����\���	�������r���w'/�.�O�o������,�u��p�O
�^M���[Д���Z<������'x����as����i�3 [}^��t�X��>�i��E�u�_�2�?⥌�w7�������e}�a� �5���#Б��.����G���D¡!Z���Mⵟt?v��ۑ����w#޽]��	?�c{�>z�E�{.���oߚ�lc��Uι�G�ô��8|�&Ë���;y����lHY�.��O&������w�3GI�Տ���?�ɏ�z�����2����o��������E>x/'r�e2��ɗ���s���٭��@y��d�WK��=ө�ޏ��d��f�a��-�y��}S}b]e��r����V�{�:�$᫗�3|6��O>��p����~��Կ�����ݏ����M����C���Y�ȶ���?u6�$��i��9-�7���]�Ha���=	_�֧z�@���:{3O�L`����[]QO��nL(Z��@���CH#��,qn
"y�%8�h3kOz�1`�7 �΍A7ڌ�f'��N��gN:9��/��)<X��H�З�	uxp�߸<?��tB�!]�}9�C�ڥ:l�+���#M%X��H3�Ա���O�����>lT����^o�2M�l��K>�^�W�w3#�d���o*�}�VWL�=�C�dQH��4 �\��O>�2�O9���9!<����է����N�C��S��8��US���Qz`+�1=t�'l0���V�=� �g/cmCj����E�:�؁ӡJ�Ы����w�<�H���m�>i��%��`<O�)�c��-<��m!�������咷v*�A���� &@ٿ^�7�am�>W�╿:�������~ҥ5-.5wE�_��O�8�<���p���x�q���ǉ3�����U�ҬN����e$���u��T��7  @ IDAT��[m�̓_̓/_�p�~X��m�h i�$+\�+/-���%��e�\��w���.���rO�{�gk�M��HG���)��_��MX�C�� ��O6-��z�C,8�`�v߫�B8򸦋w0/�8���4M:��)o���I�����*�=�+�:��k:J9�	���Ρ ���'N��#[L�f0� oO��O��f��{��mp�\x��z�W0���uk�����٪beyV��r��ħY~����4�y�ԟ�����5����l�Y9��}���Iw���E��y&e�룈#��%�LH��.��7ma�a�֮ץ�޼���z��g�Ǉ���?��w�W�_��燿�����ǇǏ?�{����0��)��G�"��שk���o)O��;y^�ա��8.��rXB�1�]�-�UvS�R����^�eo�Ē�����|t�ӑ<Q�-���{�)��gu$ß՞�W��~�+efk�z?u�ֶlẻ	���x��μё-S�âӋ|��$���A&>N��>�}�g��=u2�(9�ń}��u�z��Jxj����E�.�'�Vd���~q���{��i��v�^�E˵����B���hTC�sŇ��Aޞ��SIx�K�M�94K���b׃�48�V��.�	�8��K�2��+ޫ��2J��J����&W>{�G��ԕ���p�߼����7�lzjx:e"]>�Ni�{�nt�J���k<�e�!���/~����/.�xtXE\�Q��e������'sTܵ:��{U���(��Kw�^��wI6���q�[�B�y¦Un��`���"�=�Jk�c�0��iЕt/=a�<-��Ѥ^�%ӏ����=��*u(�$Ms<hPH���o�>�
�>�Y�6���{ �pzaǀ����i�[\2sBplC��=>:�%��L�َ�`ۯ�%mpȾ�K����q���`�Xh�k�Ȍ�Ů���[��n��ZѺ�w�"��@�Q�G�;z�ʣ0�7Y
�|���*_����q�f�hzi����s��fY��x�^��6�,�̫�<<���ꮄ8�+G��&#?�Y����3*H����>�nB��@��K�X^�m[��˽,�}Ow}�f��ng`�&E��n�<̓�����=W_'��YO�<Q���^.���`]&��\��i��MzF�e��e��[�"�f�;�`�>ƓL�d�@	��O�����[r_��#80��_�Y�&����lGQ*��N}S�q$f���M.��}-n)����٧���9�hlf��Q2��7�N��я�(��?-�����[a��N�,Ktw3@u�%�o�+��=9�=��i�P;�Q�P���?=��'?9|��-??������pg�����;�������4�"�:��w<n���d')i3Sw�}��+����n[�Oy;v)λ��95u�)�`�%�^'O�M^oͻ7�_>;<ϷC�<6tl�sz��<1��py�F9��;&w���ˣl��&���g���nٺ�k�9�6c�����e���ݏ�H����3�,�er�ٓ˯�}����N�I�&b�#K��2w2��_�h��5���6��Y�*v�
e
&�{7�%>���!H[�W������x(_~�u���HGzq
+��B���CS+lyț�p��o�
V��k��nْW���n~��lG�%�\e������ii����ASe���>}24�4��4�*��]�)��s�i:>��&����Yuz���\e/�Es>�ǋ]8yxYq�tq�i����GƆ�棞�'��?=�9θ�ի��m�<��+���ػ���A�t�~B��/^��^�x'B�[����}���m�Ó�l nՋ�V_p܄�"��J�%�<���32Z)�h����/���[�8��6[IAgO���V�4/4����*O\�Sy�u��u�ºF{�L<��Q޹p�Ѡ����W�B2��p{��0���m�e�:x��<xIZ����j���0���C�+�Vݖ������ImR��ɵdm}@s�]})��U!}��sD��jT�E�����OT�*?�w-~e��kx�a����9�\���	%:ջr�[��w�A�o����Qi����ܖ=�ȯ���W=���^��S~a:�K�4�\�A����+���L����8T4oa�}�r{"!���O��V��y{����>�
u�~mFzhG��TfO*��C>e�6��e3�n���q�wԾ-���܋����@���m�[G��w)�L�nۃ�m:�?^ۣ�ǥ�.��F�3�C�*�r�^��Y��U����{OG;[��G?�Q�G)Ü��O��?fRvy��O�(�ۇ�����?�������I�.e�:/��I��M�0|���R?�Է>���{7S��O��~��ԏ��k�_9�S�j�=�Z�g�Ux�'Kk��������H���k!��f��d�������(����a�^���/wL�z�gRw��e����G�ʖ�g/�5.��w瓜���Cr;9}��L��2�a�;w����F��(�"�T`��ۧO¿�-<3����G�Y%����}���z3��B^�cuj��m�!�Ŷ�CG0hӒ���5�h���թn�K��@����Ξ�pml��s�O��b; 	Ӱ�ذ�ߊLV��Gp�i<GWn�w�҉�?���'d�"�C�5��X}qf��I�bCKi7S����:rFx�3nd9�}(���h&�A�v� �,|��߬������5��i����������rN���W�q�CE����Mրft�5|�^�&c�	�m~'��(�+������{��u�I:g�����GV��>�l<E{�Qszk<��m���v�F��Cze�D��&���K�`\O�CV�<<��L���q�| &\yKW�9�
{Ay ��aP�.7�ֻ��>Ug:�+����Vnʏ�k��ض��˿������n��(әŎ9�[�ͥe�.u*{I[G�gp�:5O["Z�"���u�%E[TK��*�c/�~i�6H�A	��&���N��~��?���+�A���F����)��Kr�����p�R���g�4������s=f�Ϧ��@�91d�o���	�I���G�����d��+�=U���=��ˎ×�֑k�Z��H�X�G�����c������7�{��\�C�������v�(�C��XG�㤧7JSy<9����N�Y��#_�c�}�m��z�
�~��D��ה���l[���et���[��Q����8uSN�y#��B�7'e�O&ץ��~�<
���W3��>���/{�w��n�to�G�����+x6�o��ߺ���}��78ϓ�xtƧ_�}�Y�$K�02�z�p�;2\�OyN�Q��œ��K֖��%p�����&	��������Q���/϶�ց�ا:��T��%O_��ݻ���a�}�������=�i^�}��\d���8m!���3t�Ç[=��	;���k!7v��bm���O�D��gCVy&p&qU�78�9��7�����~cVi
ݫ��{y	��'��E���?�j��ë�߿�]ϟ�>�}��9�(ߡ� �f�T<|�(𯳪��Nx>^��Ӊ�LҦR�S>���{�IZ��`l���F�l�:�c����=�U���i�$��f��d�q;���5e�n\��)D���y����g�t�>��'9���W�����������d���W���Yt��_��p���2��>r�d���H��}��F��x����#�ws��û�>��_��I?�n�^&[/����f�篧.zO�=)�7ެ���#�gԧe�ճ��"��e��Q���s���j��+�����i���j�k���qp�װt�u�^���5��ec��uw���'Ce"�N�|\��'���+oq9��w0GYKw ,��[�p8��&�vT�C�F����TA�|��0}�|�f�	]��
��1��}�w҆^�ѩ�G:��nh�Ұׇl��ο��0k�JG9�\e��JGN]���V���̪��q|��������b+#|��N�U���r�|�`��
fM�~��s���n�=���i}��'W�sz�q񻲅��-.|i�'m��tnh�K���^^[pK���̤w|�h�
�n_Z6�_rgR�N**W�ꀞ���6(2��a����dMȒ��~&.�ii0D�::|x�y��뮲ܖ�fxU���Kϥ��^�+L�Ш���5�����Uޕ����naʻ��^�p��u�*C���^:�S�g ���-��k��sE��UGi\��7�,.�`�!}f��I;�4֏��4��� ��3`I�~�����z[�Tx�қWy�.�P:W�{��rx���KG����{]���.=;a�V��Qt�*#�<WY
S:�mX^�(+����mB��'S�+[�E.�����;.���NiK�����<x��]�W�}>:��ߣ��՞��n�J���s����/�-M!��|��U&����>���y^X�$d��<����/s��:��V��2fx���f�j��'^jxm��6v]v�c�:m��&�ƥ�3�A���v��n^�?|�Od��۬�_dq�V�[�w�Gi�&��3�����'�@�\�\O��c�_f[ԫI�������q�ĝao&?N�к_l�('>"yu�I����<��|�>������×�d�Gש��'�/G�$\s����F!�y�B^��S
"��B@F�U�&H1 W���x�X���^{�wV܍�*%�J)>��f=\�ɵе�>�<���08Xp��_�8�3*���õ���zz���5�e����B�V��U<F��4���|!W��V�HI[��-m'O��6n����\��������r�����f��z�OZ�B�:b��R}'?*��w�k��G���v�{9���~�N��ڵ<��0p�\�l|�&�+w/��|l���3����IE�'?���:���O�Щ{
�G�����
}y	٦��}�k���t���v�4-w�I���Zy%2��r�3������h��_�7�x���c����n��┻�:���w�u�&O�k+�����[�Ȓv��3:��	��|�����v��\q]]�<'_^��-��(?�W�ҨL�kX��P�҂�	�G�KC��-/i�mZ���!0l�w���%�e]���0#��^��L:Ȟ4}><W|u�,M��F;���!������u@J�y����W�:��5�c�����!��ڭ���'O��{�����<��;�o27}��	��G�P�>�e��Q��|�Gy��;��]�Q\q�?��^�Z\Ȗ�"9p���9p��4��oˡ��x�q|��ҫ�t}�o���VYaa����tWڢ}f����a/�^_[���M���ע��� wrt�>�����7���������yV���s���ȓ�_�]~��_Ŧk�86�8��R�e�����]�G��*cK�f�y#}���ݞV����y��E�<%������s"=���lsR���b߼�x�'o)��yR�}��9�)������c�L�^=�S��D�6����̹ۥ�g��i�1$b�	I�v�䨼������7�8��e^@�֩��|�M6B�ꦡsm�m�My/��ŵP��Zy��_�[	��BϠ&����8�U��+�>�m[�Fā�����j�,y�{���xaCr��j��`�cVɳ�@��!�Pqx�-�m}q=�n����ٻ�(�-�IX����/����v,�E����h�P�=��Xd��*ǜ�`^{G6��5�1��7_|x���u����'�*����,\i�p*�<x<��v�������~Uy�+tݴ=|z]y�-x��Fx���i�w%�a��&�t����n�kS��Y7^��m!�Wʫz	fG�ץG��+�Ґ��7���}�u����7��A������#�&���=��w� ��N���G~�B(m�����g�!n�[���d.Wz���:|q�Gӆ@~��hWZB�Y�ޥ%����!�NڑW�n�8�����K��s��G�-R˷��S���������p��� ץ_���n��5.?��0[9��Ȑ��Y���˿����˻���'8���J�*�P>��:���V8�p���g�����z"��"�6|� �����<���/q��M�.ޣז�w�ʷ�M2���N�N���[��t���o��Ŋ���X��0N�񖎎��0!��(}��iO�ޓk����U�N��[:�)�_Z]�����K�=~i���W�<���g7�7_}ux��ğ���G����=>��ӿ:|��7�O���|�U��_}���?������Zpc�S��꿧7����,6��:�`1	���	Eڹ	E^�H%���wî^��tt'�����񩌇�YTz��G�^^��e�z� g5�V7�3�����������9꾓3q@�0�'�-Z'��E"'+�e{�E&#��E}�'a����o��}��<�ޑc���FtOj�}�z�|0�`�=���"�w����kL�pZ��}��
|+H�ʢqq�0n����()�ݪ��^����Û���B���1�e��Ϣ~�R�*L�I^䚺����5 #��;ʼ]�; r�o8����-�t����xq���oKw]��[{N�U�¦�O��1�����S?��g�
-N�&���w��/�J8+�<qh��sn���������lE���x\�'��*��SVg�~�'�4*� ,lCi��S��뿕�VO~�p�nn�[�iҿ͕G��r�;�i�.����p�@��ݦOu����麮��o�H��d�=qͫ,�JO��7��ŕ޸P=5`���Q�B���a��ϵ����_�@[���w�3��1�~���|G���G�Σ�y�% dLZ�ҟ^��i~�g2��Oٷ>����-84z��^qy�V'��8ҊS����	\iF�|�^�ݙ0溲4}�[�n�Z]р3�%<��f���:��s��\u�;��Li��le����{x8�I��-��w-����óMG�u���F��`��y��5?�m�{x�]���+<\i�\W4ܓ��]�K'{�k�:�d@q�2h5��o%/��	��n/rmBA�zt���p�Ƿ/��fSN:�GS���i�'q�>�;����n�)�^�w�S:z�k��C��ⵏ4�{'���qpW��Yai�k�_ǃ����+��m��2��y�k�ϯ~���?��?>~�������'�����������4�W_��<�^f��w���óg/?���	󱎤�OmJ���b�lO��� 7��vލ����Z,�4a���'&�ܜ��I�wc����m����Ё=�`>��*���.|�$��ӛ>z�&y:��+�y���=�gF��0g��z���gr#m>p�r1�7AV,��κ��c�6�*���?Cݫw�Vy(�^ʖ,��*������>��-,�\�]���<���G�zו�!WbF1��/�(yq�|��n�&���Э7/>f�=�)J�oRѓe>�	\��#oWV\���ՙ�{�~��ʫi�i�[f�]������w�k(���ku�iH������t�;^���σC���7�7
_W���G�*����<�Q.��{&�)�~@5��8���z/C�n��Ҭ\�<Y��I���^]���{�_�
�W8�yU%�����=�OZ��0A����1!x\�T��Z�h�+|娼x7�rO�v��a���6Um�=Q�hGz�:��:SG�}&y�k?^���z--<l}W����h%8C��V�#{����皶�aNҤIGCȆ����]H.l=|ym�{�*_Å}���3�ܝ�u�z-�~Mk���U'��艻QWNit�l����tS��|��|~�>����{8�+�;L���V��������h)��m��W�ď>W&�-+uӀ�u]��q�k��/�=l�(�v��V^��~���o��n؉@���<8�''Y�JS>^��2��'�ڡ�z�,�kx�W�z-�R-Yї�;�B=���u�ɇ� ����X#���fG��o�$�u�U�����s�ծ�^wŻ���.L�꼇o~����n>:����ma�L�~��������燇��E�[���lC����rږB|<λ	�+�	��|��M�o��n����Yx��9/HD�<��i�w���V�,���A"��=i��EroI�lu��K\�ԦmQ��,NϢC�^��	�.�������^䤯{3�Y�L�y�Y���u$-�oG�� ~s�<%5���yB�9����⾳c�&>x�Y�jݏ�S�w���`��ġ�
]5����o+||�k
(J
Ub��*�x�{F�"��Q	�뚜�)��Ǧ2�|�2��D�5{K% _��<�<���O�90��CɊ��䇱7�v/��)�G��?0C+����ot���׉��f��7�?�+�ӑ�Λy�c����G�I*�1L���Ͷ#3�<gɓ=��3��$���w�N�x����mZ��5W�j����6�5�������Z��_kp��Wq�X��;�m�AZv��!}�A��~Ciu�ӵ���k�fDT�J�+۞�U��ĩ�ۛ!xn�Yv﵎S:�	�ß��0�WW���x\ɪ�(��Y0�*bD�s�I�7���C;m^��-L�n��F)8�¯n��(G`Xf�snV�C�������]d%2¬�F2�<~�Z��<���қ	GH�^�<v's|����q�U`�D�j�r�,��~�}hcy���8l������=�l�������䣿w�紶��/�^���px�,�-�X�9ɪˁ�2��p�%�r��-tp3��W����S2�z�+��R����Y7�oo���~�oq��>oz*_tfpXqi��߃'���}p�+ce&G���7��oa�rB����#=���ڪ2x�B2�,o|[�����]���K/�0�oxl<���ci��8O8�6�CJ:Z|��N�������+[uCG���OJ|q�����.�5�|6}d�E����1
�8��]�βX�p�����FÛl�����og �����8����4����|x��y���j^n6�{����=2��{9y�V�l-��O�`^�I�*wO.O������*[vv���8}m�v$(�y�I�N[VE}�4Os�8��O2a�:�I������Ӌ|�=R��əӠn߾?�e�?��컖$;�.p�;�\��$�IYZ�EZ�������\\���(������;��ߎ��Ii-���DfĎ=Ŏ1#3۪<>�,�IL&	�G��ұ-�E���r��S{����7�yk���ܩ`����!���C��7��NQ������j�'���8���5��X�S�:νmѾo�8C��kŜ�Cg�#��pkk�T]�J��@�8#S�V���Xa�_r�h�U�qR���V�	K[����q�����҄S��O��ǯ8�<6]]7~N��Z�|�i���b�D�)�)�4�����ۗG��#^��|�o���?�s����ʨ��M���|�����%+��}]��A�!n�ļp@ܞ��Dl?#G΋+��[t�p�3����#��#�!�t�ե8�_����~���pBb�?Qs-����/���p��5������9�4�����7s.za����0V������ڦ���ҋ��I��<U�r���w�K��٣�b%6�5}�hOB��-�|B�zmS\�ꍃܕ������[����3�H�q�2���C�(�8xM�pW�I|q܁(4���u�G�bC��>���F����Qi�ly(M6,�#�m�=��q�3�"�	��`@^�V)Ưsև��[y�^^����;ʩ��TN��$�s�*o���|�j��gP������Z{�4Oˉ��o�8��\=*�뽞�\�gL!4� p��v0�~e�F�>`Kyе�J��Om� �s�7������^��  |x�8�h�c ?��ѩ�#]>����s^*��׭��� ���M�=d��������Vi�%��c�l5�Wn��;��?�C������'��&� �_�Uj8��4ۆ��Wڗ���lG�Cv���:�8�a��G���q��֝E��\��Y��W�{#e����<�����^e �2�w�n�F'<�򖦳<Gq��ͫ��^eGϻ���L�>�<<�7(�����2���e���k3�k����I|�'�j��"�/�*P{�lх�עܤ��*�<������y��(�-� X���@�)0�-�⬂�w2��u��O��p򎉇�Y�W)�s��Ny�
u�+~y�7�v@���#C�i�(��]������G%�idȌ�j�B�ZB�-P�R ��<+
V��Z/�T����&����s@t��$N�/;���4<A�̛ �C�U
y7}�*�<�2�>�����&�����w'E���>�@���,�OI�=��EHL��{h�D�fWy�YpRS����!v����	��kidt]�S����;��������۩qä����� m�V}竗��z���ш���-_p'��F�Ԑ���%�zD�Љ��tR�\���X�EC�c�����I��������K�%�h7�����޵u��ƶ�����q\=�M�s�}WE>�P����'i+�>k�A�ӐN��)�\���DD�)��3x������G��9ra�ի���s�����EN��	�3~� t��-4myɫ�~�8�bi3L������B��غ=.xB��[ǋ�k�˿���F׳Al��§P���%�5֘ql�uV�n���1�6�d����v����|�ud�0��޼z��3ғ`�$��������u1s�Fs*D@:E������4�9�6">�~�G���|PltZ�$����z�8�{�Pl�W=oRfk	$�[�"�vL9�����LN�g���օ���������Z�Wާy@����V�a��7�ޥ�����+ޞk�NyD�VGt����ٔ10ȝ2}�����B� �>g>�9���E�&�-��5�Wg�w�.��o�!��̶��G�C|G�ȋ�kz�|dN�����m����2�gp��ϥ���Gƴ��Y�C���-����.�H��̢bP���x��H}�7ܤ��GŒ��ѓ�m���O��=��1����
�כ�f��]_�2��1�am��B��E����6��s/Gq�dd;2�v����s��q=Q��@3�b����kv�qb,;��.���m'|<�7��j��ůe�%��7ϐmyG���X~\��.£��j곟���7(Ng?��������͗_���eP��'>��ᔻ�x~x�ᧇO>�"w|(�?� �W�b��Z��&u�$�����mKgo����m�mƅgy �*߭�H{r6B������H����?o�:�d��G_��M�绫�׻,ܤ�o޾�� =η2��f�wi.��7#�)2=� �X��W�uk[ӣ|�$�����!����s��s���arW���ó�L&�rxw�m&!o�����c�H����P�\^<�=.��Z�81�QgRVk��&ɵ��h�O��i؊�/�q�]�����iLS��9R+B�OLl6�����/�8�ؑ�v�ř�A�c�%^^dhCR�s򏳮�8�#���Of��Q�M�����p�Gq���O+���+Cut]؟�W�zm�׼���i:liqNmqJh�A��P�
*]���0��p✿Wr/�l��eu��w��sa�;��[��Z�ۏ}�����-?�+����ƕ��Cy�+�����Ɨ�ujh�#�2����`��=�|W��c;���o$���^�%��O��FY�}�����T���z,�+Hۃ<{��VZ���PG��y������t�����!.��Sե�|��o�N*�iJ>?�i�B�����eG{�B��Bq�\�>.N�L��sq��Nㄨ�&Y�[y��8�����z�/���/�N�T���߀���P[|�#�Qq��mF�mb�Py'�칕�B�Q�$�;�y��S汜�Ǐ/������dq���7e�^�*c8@S��p�+������S.�A��.���G�tD̄Qy�ym#}jC��6�J�d�s�Bo�����/��'ɽ�L�%��Y0��䟴��wpk��z���yi�9�[��gh��䉅�'���k, ,�:�t��G��q�";��^xV��� �K(M>(=�Z��Z���N�ËK�5y0!�������˧��'#zG|+���,���l��������t���0~�A�/��d��	/<�#�5:i�z֎�MN�s�т[[:��������x�Ѥ��k5/_��-���z�H�s����?ϸ�d;�8���l3�;�$ ���I���(Jfx�IHڞg8d���epc�l{�I`�k���b�h�IC&$��\�:ot�� �W��~Y���Gп���^}���]��a��E�>�ȢiL{�	�g"..?<\<�7-|�0�g���2¿ͤi}~�����M����o_E��Ó��ٌ�Ë|���w_G��1TV._X��-�\w�!'�r�*�X�:�Ϲ��﯋WA��7�z�l�3K�@p~+�O�҇��,��O(�N���Cj<��
q!�lˉx1�t&��nN@.��苞J1�ik�Tp�{�u�^���k�������6�W|�9䊍���ơ�lq_Y]τa+�(muf�H��Oǻ�󗐘��=��f�Ŷ�y	��D��
��ܝ��럢�	A�S��߁�
؆��y�#���J8hW���yKO�dX��kPٝ��i��k����.�Wy#qLh�%�Ef��9�����G&
o2�+��8��N���w.���,i-��!(��]��?��:�]�/_V_��!z`/ϊ�������5;�S7�J��^֞�)O82F�!𚎷�`��b���e��S�����&mV�Cw^818���U����4rO����>͹6cڝ��/��7��L镦��ս!���FcE��_qKfq��4oy>��twmڮ$Ӕˢ�l��Y���qwil�Hkz�ˇg�v����7	�;��ˏ��'�ҜA�ʅ��T~Bi{^ʰ��vˉ*K�7��]�ݴa:�g��Fe���W6:㝪��탍3`���L+�U{}�lԎ,t"�RM�;(������0�ȃy`�^�jU�7�hxk�¿�V��������;T�Agi`��"r@:�+[�U�`����䥇�.�r	��c���[y�o�J�[ڒm�RY�?��!�j,�8�u���=t�u�BZy����ʉ�8���oZ��o{y�;���s.>�`���:�cH�Ό�����2�/"2hݶ�E�gY�� rjNd\�� m����ݮ&�r9/T�^7��_�����<���E���]���p��=�s���~1/ÙmJ�=i3�.�_px��㼦�2��]�B���Tİ�D���ĩ�)S:����g���}Kq�LL�݇w�����qL���w$�\I���@�d�s\��}�������U����rv��s������*w�rg�ݛ����2��%��:����9|���×�yN$߰ȝ������Y�\��)Y\�|1:�u����p��O���?u�S8߈�\����O�BM�T�:X�5Ѐ�9��]�;�UN�z*��T���b�1KGk����ek�����5t�l3`������K����&���F><+��jk�%ǽ��G��-]�%?9�~��UvtZ���(����!���3x[�<0s��k@� nX�\R%��5��[>����<,��%����ɹx׀���_�څmz��tмʮo�@Mzq�0��v�7�����Wg]SΛ���	DN�o��r��|r���yhn�n�B�Ȳ��/����u`�n�����g��ۮ���/�.��p��=]��[~Mk(�n�����M��w��O���K^м�e"�S{]<�:_�Kߧ�;8I&G�{^zk������M=Pb�E�颗�� �h����F���v^�/�q�ܦ�߷���x��랣Q����G�I��J������^���Jr�pYP���%�J���-ֹ|�:o�}�2(��?���W��e|N�&�NB�T7����ߡ��.?&c�lt��p?���G[�˼m>=܉�n�6Y��{�29*�}⤰�eC9�_���CdO'��Bq�����&���f|'L�8w�e������������!_q���ԯ��2�*�������	:�=n���Sg��59�OqKC8���|l�|z�=���(�$K��^#j�P����{�k��x��Q�x�[����[�֐���o��r �����p��|��4[�}�v��%���\g@�nt|����c\���_�/����Q�m0xN�T������O��8ILڲe�%�Z��xz#ңG7��N�>���蹶�<�j��|U�*�<�lo�ק&L�p��g�2��\�|k,���X���4��f9�L���Ͷ�����ΧY��o��S�([�.m7ʛ�B!��͝��y��i�?��|�ۤ�N�c/b��<�m�Ӷ�4cTx�x�|�u>ꗯ�_�c�lk�.߿�.w#��1�}���ѳܕ�����i�%�Tkm«�?��~=�����P�C�4����K��6�hڜlxp����Vڌ�t8fo*����~8��ϟ���m�����Y��[Yb`ǒi�/�^�x+���V2!��@�H��M{���D~ �>Hy�9��\�2��[�I5��l=�x�7� ���)U��!֝����'��C3IG��s�|�g��дz��{|{@T�M_ע���#�����������q{���M�vda'��ɧ��9c��~��W��S�����NP���6���.@��\��2�kd+H]��2�VL�b�#��f�S�._�k|%�u��d�<�aj�ڥ�ip�O���A~�l�/c�4Hȋf�V������Z�x#���7_*-j?��s7,8�ax���.�{�x�p��:�EW=�ǡ\�����ǾB ���'��d�6�9��[�#N���t�hRt�s/�p>v
�NXu�:�Bi��n�n�Cw;�^����yu�ǛW|
�y6���Ã��(��y�rх��p��Q�͎�J��z(qBm4����N�JKܑ��SB.=h?����v��Ix��p�{̻ɋ�_P�\w@��dy�;p�kd�h@t�����QW��<�|2�걕R[-g����p@i�E~F�����l�#ڂ���������y�t��&�&{��j;��W�M�Io�3����k���2���w�FY�>��Y�A�Ђ`ǡ�Ub�ٰ��T�����+�v��I_^�w���x���/Y6��lsIy{�o_7�Υ��s��ܫ�ص8�|�K�9�g����]�_dbD���m�/���st�S�K�� Z�����4�h���ٳ��i�z�C��SP>>v$�q|��e���������?�'�>|r���O<�(~O�ܩ�����z����7w�!���.��J�M���Iʸ�<c���,VĄK��u�x��[��*s�Nb�G�Z5ߵ0�Ǘr�s�4w��}�IM��位�����*۪e��mMW'o3M;B�W� ]|�ￎ�F�����G��;�"���C&+)�Ù;.�@yVd�Gʫ�N�Mj�+����G��	w�k�kÔ&�O� ��<����Qn��᎓׵�x
��Ax�7���_�ռ���:�?�V�BL��#0����$4��;[^��ʲL��Z��w*y�Γ�l�'�����΀���-�+m�X��-�k��8\q�|�ÓV(m�#96��H�|�L02%�׀�4}�}�6��%�1+�yf�����*�^�a���ht���G��|p�omFє�&�r ���,?�o�^�[u�[��`=��u2��{"��C��G�C�'2���n����f� K:iy�[���Ӹ�\���c��v]ZItJ��|��K���c��4�M>�m�:�@��t����4����]4��#���I2J�u�����"+��=��s��Ζ$GgdY�:{�=������s��|ߟ�����������t�h=����Y�������C,' �U}NУ"w7?�0�x?a�=���]�-���r0x�����w���� � ��I\�)�(�윱�m4H0�0�q�m�e|��&~�.`��y�)]�Gd��|����Dd�=MA��M#�#�z%��qF���+S2�nﺺ�f?�\��A�=,�o�HrC�R-<��{���4n�]p���ݣ"���Yc̡a��[뽱!�"H�F,t�/A��\�#�y0���(PU���i�g��4$]��|W�'���J��Տ���KR��t؀-�%]vBj�Vb�xW!�2&ͤ'�N�>��}y�w���]���o->;"��Pɽ+_$1f�G~\���[ϣ�e48���#�bj0+Y��s͈����m� ���A��R���]��7��mW�i�KE�0!��da�4�ѕ�{%�j���4�ȵ���7��]�E�m���p5������k8nׇA��� K�HdsuԄ��	G��$�-#䫪�&�ugd�@��ֈ|�i���h���h�9���N�
���oݖ��&���jv\ł}�����<m�s^�G�g��$��X7\���]��G;lu{)��x��l|��k�] �ԾY�d��xa����~~G���2�����W����fm��O��Я�5������Ј�o�����k�?����νl_T
j���[œ�scd�gb�:�j�4#��alk$�ܚh�WL���v�[Ț��^�.�t�C�!#|ƷT��$�p^|��5�v]z��˂0�IѲ���&�5!��j}�u_��گ��g;�����<0+��!��w��M���*���7�J�}�#�ӱ�̫��Ъ���Cf�M�ִ��u���b:���#�_ך���h�J����B�Lxs��#.�c��R6E�K�k���̱3�4��@�7�W;�����lX�-�ύg�\���s���BJ4�c.� �#�t��=h�f��ck�^��ԟ�]���+d.7�?����zY��&?��]��V������z>tes;�t�D7�����K��Ov��Մ�rE�1e�/�}�Z"�+�۳����	ۛ&�?�8���<]bv��\bp�N��vy5b���uͥ�d�v3�����y��(`��g���/�3�/6$m������h���DgFM��wmHϮ�M4��: ��&u�A���BE�bo�Ā܅=P������{W� �1�z9�Is,�qD� �Z:��f���<,|�g����v m����
�v��f�����h�$<�֗�c����Vc �9M�Q9�[��|,#�ϰj ��p��g;$��Eń��(���a����+T��Z�{~mo:�q&�Uɩ�}"xV��`�0�
Qc&dU�E��|�w
6����f{�%*IIR�a�-6��ur���5����+�E킂���孳���`Z�n�ݾ�g[���u_�D��J�R7s-Ѣy���a�tP��Ԋz�*��9�iR��>Q��Ȭ(��n6׌5��W�K�����N�y��4?��Y5�������mY�o�[vߤ9YA �uWH+;�Q���;XcO��B?7�(�^�_��;@�] ����sb2Xb���p�j�؀\�AX���\��}Œ����=a�� ����Z�'�TJ����<k�/_h��2XD*ѹ'�5V���Ujw��r��vf�8��udS�?�NUT�U���Z�#jJ�?DDb��IVw���
��a5�:P�̂�n��ĪX�D����i;��'f���@Ƀ�?�"b:�J�� �Ļ9�r��xd��m.h����z��Ơ�� Z��7�w��:���K�a�ɖ%*ۼ�C�����Ww,"��s�0���7�l,`
 �,��*�p2Nj���p�Wq_��-�nZ�/@�`��lu��0e�R�]��e���;����]vD�����R��6:\.V��1%k#t�.k�����h.��A1Ƣ	���w�J�T��j�����yO�//�r�|�,9��sޙ3���˄!�屎4��UyR�izj}�~��I0�{�A��%��%<�)�@��[�n�n�ZA��o��xw[҂E�|�����>���Mf 3���&U+�d9&"0y,0��@+�I���{����|l�E&��� ���St1c�>c��S�X�+�Pm�ҪNf�f�R��������"	�2`�	J-���	D�Zo�n�����6v��s��e��ǡc�X�0���Ɉ�Ɖ�!l��0���%I�7�Fq��W?Kk����B��ŁvjmRr 34V)k���b|�&wϗ�\nA�'Z�N	V�x�����k>�%����k�Š����!
�f>n߅��q�f�m�ü��7c��G�z؆w}���w�;�J|�֙�:�L��"�b�OF�\H�$ؾ����^|w��G9��,�+Kخp2��7l*qϚ�1��O ���\Ŏ�[ ؙv~[�Jl�he��%h��E�EEФ�Z�+��:C����P���1Ka��U����Y�����Ih|T�uZ�#dr%P��@�(�����*Ŝy�Ǽ�p�������l�y��D��@�Ώ��8��Y�퓚{�t��_���gR-�@7lw�]c�����g���m�{]Ɣ��f��{E�|�8�;n�� ������A����KqCh����rץ�v^f��Rݗ��`}��so��U74f�=��{'�A���hn�%B�m? �����#k
����ƒ�wC�=}{&�B��w�JX@W�� �=#��u��L�]��'�@8@���G[ݠ��%_��/���k��9�<2j��r���C���/�SR�g���W�qM;Ο�^���4��P�_�@�S_ܳ?��~6��퍝�7�"q�X���m����,)9���d���J'������3�0Y3�Xm����4��A�Iq�s��j\'M�[Q�'g�ű�C�\m����$I�K���p�� �k,E4_i��Ϣ���V���x��FӔr�	����N���ڔ�_J�/([#��TNqu�躨����,������G���iߞn�o|,O����A�/ �;*91��ma!�nֺwS��Pp�'�A������S3��	#r�[FX�8��h@��%�,���?D��X���i���t�i�S{��Y��R���:9�䱬y_�P����:��L���[��ksd�XkQ��=��Ix�n��*�i��jd̘����������ru[�=� z�����a�)�"W�&�
M�>Wf��Y�����kk1�_���H�,p*��L8S��{`������m[���d�BG^(t�U1)$R�w!���,�������N�G�3m�5�/]n8)��9��t�ҕ8�
!�\�k����{�j[����^��a�|�
�7ؤI�xs/��|쒭A�~M��̦I!^��Tژ�>���O��0e5m�ߔ�\?>��sݎ�r���Ҁ�1��C����I;X��>ᗟ�2i�g<wOȁ��2����nY����x�2�y9��B$��ME1��t��z6
�/^r��/_5}cV0:-Z
ʞ��]+��4������3'7�DI���;� 2�r��z/�]�d5���ܟ4�@��e;�q�K.�0�S����|�"I���^ؗ����^߰�Hy�qP�<�GB�7�l�	�OFw�9]˹
���V��Jdj��6c6��%K��������(lf�|-4�~6T��x�<�ɕ��xG����<�XH3	�K@\�r����1����]���4�3of�����aH������).��i���?�ck't=�<%���+xi1�)e�-q���V*����1�;������y�� ���({7�qc�����Π�;�eo/lV��뽨ۥ�c�n%lv�,�*�El_n�\^`ůHK��8�l͓i7O�0���C�[O-��Y��fr�3��[�d�R ȝ��ώ��p#,�n����h��%���p���������*ӹv��ocX��T,:b_�B���QDL�	5��v�w*n��I�r��.f�3,X�
p�u��ϕQ.����b������z���-�}���9�}�8�����p��,o@@M�
�e����h��r#��ݷ\������*��ez<���Jc�B4�L�N[�M.��\-=��
\�}e|�EGyS���p�E�6�=D:h|(u(l�&��R]�_�����,9�W>b��0qR1���>���ـ��%4���
A-0���u���8�g)��2�B#��<�,����qD��T|�=N�}��~��t����^��b�x����;�OҜ������65!0VM�_F�;EM�g��q�Y��-�y^kX�m%�s͐�A_;uD� �/8^�1W>}�f8SOB���gẞ��{~�����G9����!����fҳTz�:Ȯ_A�ׇlã�A�i^hާIG�45�rV��#�5��wӆH�Yt���Z���;�T����3I]mW�l�դOx���X�f&���������w�n,[У���sҽ�i>�LQ?/c�:7SV��,*o��@�s�I���X{�@�*;'���l���NaTEv�������#�$�:�7��l�;�H�+�<�3�[����9�gß��C6�[���>��Ր�[@�<�m������ݏ哢���d�nE��V�rL���v���w5�w!9�p��]6� �����|�57^_�G/3O5� u�n/cIRَ�ϊiXk�~�ur24&}�lM��t�@�0��!�'/������.Mug����F+(��0}��j�ay9g��z�q(�y�46]�^S`���񛨀���&>���ј�|�&uu�Gr?2���N��a���q��p�E����
�{��#�P�����EG�6�[k���ɔ�;����}E���%��qhÙ���t�� g�Ə�v�'��Ųmx�o:�u �t�`�X N�Nv"��9V��u�h_+�͛�s}5������ˁ��s�,0u�<����n$052<���B�Y���8g�R��p�����@TD�A���auc�y׫�#0�j����c,ؑ.������<��a˥�����|U�57Y�ˬru��r�:�;�}�m+�Ќ-�Q���ɽU,Ļ���?�g
�v����>2œ�d!��<�>�G��n�N��~��a5H��4��k8���B�*�3ԀK�i9�w-n��D�^������8�Ka�ltC$��7�����b��{X�[t1����jw7����?��$c��<-b���T��p\鍍��n<+R��%�[�:�r�{<Y�S(`�����o_L�~���![�8~㦥�RqK�ű���s�� ������r���5х��
�3Ŋ�8�͎@L�C�э؊\ֈ��+�+�TxMߛX��r|Vxw��0Ud@*<�l��jd�n�q����#=�"(?غ$�_��9�VXd��Y��9���;0_Ga3<cH�|���5��4��J/X�ψ~hu��P?�|2<����̬Uh�{{��k��6鑰6PJO���m��Q�3)ݬ'$^�&�H~"Q����4�>�|��Q�++U�\{
��&�b�?�C�h��J�RIl���}�]F-G���<\1+[@P�z� 0��/rR���Ao���r���`ڵ))���S��|0���/�¤�B� ��>������WNtO0�MS�+����T�n��Ր@��%�Q_s�� ��{'@q�h9?G!PU��>�U�Rˢ��E���j4���Ѯ��XZzP�M�Ԃ,,�}�����<��<�k����x��Y(i�'�2�fP���m�ZR���W�5d�%�ԉ�5@5�4x�fIЇ6R�dɀޙ��8;��d�0[.@�q!��~��P�{5��������O_:&�	t��Ǿ��t��﹎ ��3�����X��WWv�5��:����BnHP�urA�{��|���n��S��*7!5E*�Ζ�q�S렞�s��e]�ۧ���1�&��܋�j�}�q%v�^�?���9�6��w�
�m��4-��e@p{$ �ߣR_��LHT�T��7=��g�q�
����a9MJ��o�I���XA 2����9�Zn%Y
������Ma�@��֤E^�rg�EK�~b�D�%��9Ŏu�����̿�Ws����LJ�uZ�i������ߜ��P���]#�?R���W�PW �E@z��x��9�|�.�f)��+H��6u_<�,�+X�3�ʿ-��-�%}�pw�������GW�i�Dp+�/qO�K&�e�/���V�a�0�e�Lw����2l�-���Z�����
�׸EOQ�ѵ�i�*v��I6#j{�_��:�2`A^����B0�0�����`ȅ���b6!Y�䓨������y#��3/3N<��z#t��,�רY"�Q�kf&ʝ�Ƿ�l���.�a�G}�͡C���?�z�M',���.J��$٤&�O'�>u� �{���o��-|��LJ�U�� �_���?'�E8�;V����-!�W� ��q`�۲��j?I��Lu��w���BA��n�GG<���~.�_Y��o�}�wvr�S��y#9%�Z�Ix��4xU��PU6�0�s��#c]��k�O��}�v���m�h��*q�Ҽ��I�z���M�3I�,i�0���w'�4s9�Uܺ݃�Z�����;_�Rb���ߦK]��7y��}���27όQʥ�fx�����}㗃r�<r̉=���ѷyGe�I��0���xነEc�'7p�+q>apc��R���sֹ�Q@8lVNe�������O�'��!x������1������l޴VÂ~��נ���w���s�I%�۩*��hUȢ}�O�����qy2�����Y��7͛����c��9�o͎<��XZ3�,,��ִ�=��'Kv�F��K�n�-�9ߦN[��H�.Pr�5�{����B0f�̨w
l{������4�y����V࣓�LɄ�"�x�X��N���[�yR�8`�f��y@U��(o)q�J�Qn}u��V��vX�u�C��0��5��S�Mb�c�J��_��I'�-��Jd+*������(�M���z� �z[g��D�jP�w��@գ�t,���XhN�Ȳ���{:̋#��?Ē��՝o���;���6U_k|Ɛ�c�g5��`�0&OV]?���O�8F�#&!d#�f�����J�T��	� �����y5�u��[�%U^6���k�|,~��fR`�S��	.��'sXAՂ���љ]2��8,��������.�i�{�E2/p*����"P	W�ʙ�ζ*̻��]n`�n9�WU�+n|9��|�=2�B�*nbz�r���[�{�>x�}'�ң�6�a]��Ù�v�޺�Uيp��.5I�!��A���W���fQ�N�·%�=�����_r�^ݝd7�Il����Ӻ��я�1�o�����՛g�1S�ر	X�qi�"��ז��СW�vC���t��ئcz��������m��*b���e^��q�_���3�>	�/o����y���Ԝ��Q�!=̺Vna�����Xka�Uv�%���O��u�/�x���d1�H��Xb�������T:�'R(��[
�i�����g*�����k����~��W$���c��-���SZs�{�]ܵ����K��ZH��i�������<FR����<��]�83�z0���W��^�L*u��[[d�X�PN�{��bItA�u�O���tkxK�n/�E�ת�E����q���3���3�bE�U0��AB�k	t�~���!��G�qZV�N�l�T�#����PV#�  �!�g��D]�L�o���^dZ.i9�{�_�Ӱ42��o�0��t)1]X4�4�m�8(�0$��b$�2��i�W��85:׭}�6%��im0?�������2��a4���Rfz��0A՝U�q�n���y��ed�����-��w�n`p� �T<��ΗP�Z�&F��Wl��+%�mβS~9G��B�H����]�%��%v)R��
���Ic7S}����I�� �ٍ��6fCeִ.8|'�덌�I�[�A���j;s<�4�BKaߘQ��t�Eϱ_�x>?���[��&�n�>k���xƥ��UL��v]�ȏ�䠧Zl?��y;ȫ���?g�S\����j��N*�bB��%lL��TEy�H�2t�h�4�ߵ��:�ཱུ��<;ݽi�@� %�����)k�}���J���r�m�}ك#������t��M�u.�9�z%��GH���}�?>���m�Pv,*_#��'�$�Q�i�4�`[$�v?��W�26!G�]�zg4�"�L������t`�ތ������U��-��?ޙ>���~)���J@^��/d"y*����M?_�m�eF�n�\O�2��%}�7��I���r`d����+�ֿGi�wR�#����5��߆v��C�����v�E^LG�ɖ��1jSݥ��j�D�rwX���j���LV�9؟0����4'�����$�����T�a�;�,h�����x���}�R>��MjMk:������ ��`s?�#d���>��V�+b%��K��ǌ�u�{��~��P��d�k��Opv�J���j�pp3L����hK3F=�ؘo`(�}��-�o�s��,56'A�B
�D^B	���g#��J�f#N~����7���[��#��v�UeZ��7O����G�^&"p��������+y�+�䱣,+ro���FH�a��+K��k�T��:�?&�J_��z�$4����j\<V j�tɐ]w����e�ݙ�/{�=�B����gUٽVF�It�2Cz;#��R��6a����b/�ѤѲ����Bwe�׳�'(���ث x`���a[ci^$���P�׻�1/���t�_�F$��O1�u٬�so%?�u�����^%�l߂�`/��6
G|
%j�>��y�SN��j�K�G�Ѵ&��򥤙8<�@l谄�PAA��S(�^�';�R��կ{˒�̕�𠓧�0�i㼋`{����B��m,�����h�ۮ�����s�;��� ��xW��><�Z�J�S���_��/�:�W���筤�XX[�u#@Qͥ�x>���^N��:�h��9X�~��T~�½7Y�	'a��5lf��~�?@A��g_�U�0��・����?%7���]Vl���g<D�g s����K$���7^��h{�]2��Պm+j�fyDU�P�
��]�����4-�6��" 0o�cAc��L�O{+R��'�XErmo��R�e]�*Y]�8�N��	�.�*k�j~iRY�_��uj	WH�/��S@kVOџ��tֽ)�;3/\O�hi/e�/���M�Xv�݇ǀ�v����`������+<���rl��
�=�.`�f!.�ցRQ�>��lĎ��Bo%��.���C�3W9���b�Sk��)�i�|�����S)Yf5d@��Vt´��/���2?�������/�=���/��|�d�Q�au�_>k��A��҅�i��z
�;d�XX Di���}�,�z�ÿ�`��w��˓mL���L �}�ɲ7?����,���DxFǲ�{�9�`j����w]9�˖�W�\ܻ ���&K��%��|l5����1A��w%�~[���2U�OUk�m������14�5��\����ɧc3K8?K�e:�ϫ�=�l��m���~������U���m���4����y+�=y�?��^�"i��-��/��u;���Y��&:
��s�J���.���u�0���۵C8����P-�i0�%L<�����W�������Ilgo��*w��&�e������!ý%�<E�������ʸ�k���0��1�y�X�t�tKR���0)���c!�c����B��F����Xo8wy+�&K�Q��JL1�t4������f�D�`���5��~��4Y3n��.��Ƒ���bn��=�ƘΗ�ܲ ��t�g?��;7�6��{��
5�OR7�^׶	b���cw���[7�l4Y� ���JO�e�}1	��zC�Q�LFiQt�\K�0Ϧ��|�l����WzYzW��Eu���}ԩNdv|br o��'��J�JА�׿���ә�������a��a��Ls�9`���T� ��5$�Cl@_t��T��}��9F�����n~L�>�+{E7�[�~���X��s�+�Z�:om>��PTe`����U��v	�D�Ĩ1�G��R�������Bl���`��W����/�4 �&~9!Ygam�k[��]�6GDԹ�=%K�{�+vu!6�/>=����F^[�1{��B���Q���P]bg�恩V��
��\Y�hdN�$�(A���n�� �|�I�>|2ʔQ���y���������t�G4~����<w��(��uy_�����E�� ����{�t9(�,.�E�f���E*}�27�J6C9����S�|
���v��k�>����d��5}\~�x�t6���ntE�XZo���m�:%n���"��,��Г�Il8��RX�+��WS�?8ܑPNW�Lk!�.�W��|�P�0�R�k!?DTr��������O�]��K���Q)S"�����9=��!�X�K�~e�GE��s&Ͼ/ �o:��1�_.��>��JL�gO�{.�1��Y�t䗐T�� A4�A�-�{�f�3ۡ��<@�?Oy V��W�����-�@�М�H�{��*N;oX�2�/��M�I�^{B|�K��ɾ%ܴ������(�#�8iq��x2�2m��o_T>L�>r�.����CC0]����>0o�Fz�Y�9�`�%b��
�N���H21�����T#�Ƃ�%�g�d(�ܩ�9@����
���t����m�՛�j��
�UՖB��x|)�߼�;��R�%m4��6�������P��ȇ�mtaPit9X`�����Towyz-���@E"[��<��`Նy�K���b�IȚ�����:�?��Bg��F���H����O�R�˝tg|�n�&��cvʓ�,��ܥڵ7,�~?E�AC?���c�����`��On��pGB�]��gt%�X �7��i��S�[�4�ȠcG�if��g\�\-��_K@g�8k=KҒ����I��i�Ә�+s��K���se{ǎ�<׉�m��
��d�ԴkN�t`f��L>>���თf;�)qm�h�����'ޫ�@3J~��s��,��e���̨UJz-r�E�ɬ��ӻk��}?�N����o��.�^�O��ʎz)�LX5�	�M�f����{��`���O����+*Ey��"��vE��H� �<^����(5��n�YH�P<E(,���D��;1��?��:�������Ԋ'��/[�6�h��kV����an��56�5��_x�lҧ����Ϳ��E�B�R�<�8�&Q�G[���~��\���C���
"i�o�ٹ�D���`��=�������	B{�Zᅮ�G7�^ͥdӫ�ㅃ�ƨ,�S�[G^n�)I�Ӓ����YK�\qb¯����[ Y��T�M�Ӝ7'<6{��N�5�����;s�2m(�B�.g���JZ�k������E��M��j�d���G�5�(r� �WIo�sl�;��[�ةSb9%��%(U,}h�vZ�t����KWb���R�^�|a�b|�G�Y0�xOK��<AHQ���@�1�H�G��r�1Dhv�IO�n���4�����t�)2[�	��C�[��댡�Hw��(h�x�g��S`�������"t�1D�e�|<;�c��ͷp�$��XSou!�����_�	�%�Os��H�+V>�`��Y�Q�t�.�Oܾ�?!a��I�,����w�a�'�e���J.C��YϙX?܌��Lv>ݜ&6�X���~N��5��u(�[w��^��W�����س��n������_.<�4iYDE�nI�ȇi2K���r8P�:�q�	l����M��C�@��m��b�)�M�敷��V��`q�\��8��GJ����w$�,nܪ6��!���=x~�0px�x�䖱q�ו��L�~�-�2��K�V�#� �iLï�+uN�[hS�5�j��S[&j��g�#��,�V�tV�S��׸����A�Ȋ+p��A���jH9�(�~�\����*Y7�:X��Z�ϪN_�7#�[�f+�κ:��.;ɕ�1����_�쀯���W�� ̭I/�6k��(K��W��~���:)����� c�&7����L�k��'�`8��LӶ���;�e��7�d�wen��t>'���4!�w�E���B�E�
�@Kg�Z��Erw��!��$�UTḀ @����js�파�.�]�+�h�T�;ֿ��^�&�N�x�$x��P�Z�S�I��_$��L�7�0��s 2�u�If��"eD�N�bX�I�#q%��?1�ל��`�.��.��b�#�b{4�ɱf�k6�Bf'��G!��
ʙ�|L��F����+N�(W�=���'�0O9�а9��bTE�s��_������1�pj1gC/�:r�-0�C�'����:b/�'���K�����v���h]K�9�9���[�Q���Jܮ�̆���O`Q�	A�6X��������乌�Y*����Z����#
�t���'\<
fIm>�=�ܪZ�=x�#� ߝ�Z]ܔ�1�2S^�\��ʎ~���ق.�+� KkjK�o�"�PR��-� ��%RZ9�FcKGrz�;���RD&�\k8��g'p�`�:�N�^�aE" ���=��p�O��C2xhgN5�G7*
mQ,��ng8�� �S�����Y����R����o����M���f��`/�w��(%�p���e���
��pLIn^#yy_w`,޶ҩ�{P�6A7�+7;+e��r� yk��T���~`�-�8~]�l���f�8.1�8T�e�ȳّ��.ۘ�����9����!��k$��{�v�+�
�ʧ���&-WgW	%v���C�paF����9g�A��x�=(j���I|`�bW^5�Ti����'\�̇Hʠ������/��?��ꠃ��M�%����14`E�3�SV�L��br�([���NA��8姈�"��7�24�G�_��5�.�_�y����:l�����ۣS�����2!#|�$����欋��X+��x�N#dœ��釯��T�[�� �B;�2?gPgm��ɔ+����Q��@��dC�4Wr4O]����7"'O� M� ��p�M��3��R�J<��Wygo�x��b��V��B��سV	
�[�5K��fO34��].ʡW�gd_V��;�)9���0dM\�~�i������-^�'��܋~�>^��jA����F|u�	�k���'����Q=c�x�LWC��r�u-�Q8O�����Ч�p*����7���s�w�6!��ֳ��bFǻo ����Ds��.��й����ይ�Ys�&w��s�lJ]Y�4�dz�+�S�y�Ǹqn���Zo���H���<�#�VsN�Sօ��P�'��m�̗��xԭb��;���?d�CV^��7�/#�-��䍮u����"J�W��N}ˌ)�%��+-�f��N6T}ܛ�Kh=`���6�r>.�uC���k�&�b(�F3�!ͬ��,NNGX�YA�_�jX {��Z|�w�j3�f>���9�0�3���;n��ݜN4ޛAZ����Eb S]�[%��V_-D$���R��$��v��3C	wK<��{yv�~��,������Q�[�WK�/b��b|ϵB�����N�o>4�⅝_�M���UTx�z�(��y�d�7mQ��p�O�sQ�4)up�Vamq��xp`�i�Ә�۔z[��ز� ���ˣ��{^����tV�fjz�}1�㯣]S<s�+�s�,�G�_�ri�:j�mY��-	��n�X�lH�=����ǂG+IQE#˳s��Yp
��rZC�9�=���z~++��q�Yi�pW���ȸ��<V���yz�V=x�h�%nfT�φ&�̪w�k�Sw��uAn�Ҫ��x��5:�WR)�߭���%�K���
v�fix��3��A(��5X,���m��5�o5�v��yP	y��k�"X�i=7ꀕ�ߩHuKY�ʗ����TM�k억�C�����>h�i|��%8��5Ԡ'jJ=�8��R,ϻ�f"��QՄ��e�������
�O�f�j%��w�ϓ���!������W�QC�j��vƘ|�U8�J��	=>SȢ=y[^��R�
\� >��?��7Z8j�t�{�7���#go6��R�w|6��k8�Q�X8�dQ��-o��Β�Eֲ�
��7��S�1|���v����%|�B)���8��H���Ys ��t���[��$@��_=q�i_nԻq����#5cʕ�L�*���:�&fP#���zI8�����=�aۦ}��Ro�&{����mw�Sͣ�{������I�.i��٨-����IŦvC{�x��9���������<_f�N�\��z`t�>Pbh�ηwT����:��{\_�PK�l6�{�s�	���
�yB<�[?��S�d���<�Q*��p<�#����n�����2��9}m+5�5�����R���8+�8�l���s�V�)���~��0����"B$��l�{�_A;�H�w�x��p]��3�SHy���V��g�[y�"��w���g���ߢ.Ccl��8�8ω��\���J�cֺ�_�:�<yL��{U���.b�ư����j�(G��T��d�	]}�E��mڽ�#o�:�X����EOۑ��N��C%���(s�MJW8��A�������O+�Qg;��mQ���5�����	:��(���1��rH��Z�	����2��{�,2�AasQVGz��'�s�Ҷ��%Ӭ�/�9U�؁�����ǟ/��F�
�ħŎg^�|ko��D{_�0��~Y�^�`�@��t*򵄷C��;:��>0��@< ;η>I������ܱY�=���X�ha܅����Ft�^IK������M���q��Ĺ�h4j��`�j���*�F���d*6;n�X]�-��v,;�~�F 
��[���8ܫ�J�>˰1F�U8r�-��e�����-v�$8�fZiq�6��ԏ�+oEI���!15���(R$V఩��*l���#��U)wAaN��h�O��zǾB���-�O��7=�
�f�M��%�uu��ȼ_�"������hQ��x�3w{V{����Eu1]��,��痛����	K��@���Cu���֍��{w/��vA���T���w��Q��ǟB4��2�@����TYs�KÞb됆j��p���۔��঻gYFC�8������/�/��M��`��&{����t�%���=�o�u-1{�8����Y�%�dg�Z����5K�8l�������W+�,H<#���#MA_�.u��*��8|�0�g,*�>={�lM����,�A�]Ⳙ�\8#�r��C7�%H]��ܿ�����m�����#S�~;iǄ��'v�M%���+�cϹ�`�N��~o����ǋ��s���A^~؍�Ww���g�V#�4a��g���@��8~zu~���,gQ����Yռ�p���Q��s�(��W����������2ˇ=����Eٙ��Ȗ껟G��l��4��OoX�Wg'�����72(����,m:��W�����B�Fդtg�'�gʢ��(�Yy�{�~k��7k����ڱj��1��;/��g�(
e\Oeg��h��}�a]�<0꺟Nsѣ�և���B\<��-V�^*$�=�*�^��ۂ��N���`��.Cc�َ�]LC���G���Js�"PP�U���<	�Y?b���d�E�S�*�!TQ�ζ9��,���������W&�n��H���װ$��n�8,�u�t�g���G���;��ܭ�3�W	S$-��&!$�u�%����~k��¶��J}�CEA�)-����R*�--�lCD@D��)�!����=�XPc�����������8i�L�_'�.����x������[��^S��*U��湳��{%���P'�y�.��C�!31X�ַ�{�Uj��/����H7����/d�V��- _���vNW��V�e�y��3��5C�^[��G�����}'��F'Vͮ ~�O�'�ᆧ�!��6A�|���#��	��e�p�~J5I����,�u]ܟƍ&-����2�6�6"�yg���)���3��|����M�qTq�d�!Q�"rW��K9���YV9����u*�S�=Μ�_}�r�[�YZ��L���j�� �K$w��cP-�r�O�:��Q���0��`�����t��,����o�G;��з7�_�n���DJ��-v�r����SjTEiO����x�nN��}\d�
�4�2�em���A���.
B,\��=���Ž �e�-u�v��B@�ho���M���x�
~[qq"�X�ݩ�A۳c����Wlr ��z�[�9����&zt"/1o<��ъ<��-JL��������FS�ןB�z��CT&�P�$���A(�"]����F�o��+KЍ�F�%�����ß�w���`����)E�8�I��N6y�`��<���Bk��E��x�ຶ_%������#�^#JgH/��
Wa_Һ�5񽠟�Ϧ/6�6z_=�;� i� ����<�xئJ�$z�x������P�̂�M�f�(!�S�e�һH�=�'�FF6�i����!<�AY�CO�2�5�5}��״r+�l!�{y�6J�Z������c?V{�)ZPj���FU�&�Z�axڨ��Bu4I謨��n�?��kiȆ5R��)b~k���l��Oe~Z���;Qx�M9gհ��;��l���i�W{����f�י�d�߉��/zr�<˨^��m�Hg<���~:�mB��/zl�_����3�UD꒰�=b%5�J���8D�㰌�����ƣȾh�_٧u�H> ݯU�c��D_a�/��e���ѠPi{��p�nT�L������X$�Ě���Y��mIO�vDV��r���pu��,>���.c����$NK��[���a//�@�t֜2�L)���S�N~ByT����g���Q;�e�OQS�M�R���Y5�<��(vtj�,X�.#�Gt��I���2Ցu�P�(
�tK\���ij�6��츓�����;�.��x�C�U��5T���>IJq��U������t}d_}`�����?�����z�{��A�	��|��ᶔÿ^1$�în<��φ�	3��^��� Օ �C�GZ����Ziʀ��M���A3�����X���'��C�-������9X�_ɍ�L9���ʻb�}dn=����R7	b�y�o���ݡ��7ߌzo ���Ɏ^�d�H1�+�-yeB%RDt��7,2�-��V#<[��3�F�,����[Hz)�a���f�Sl��-�����ׄ�8���y �RGjH�&������٢��Jyiob���nv�V��ߞoL��y�d�[�	;��W�`>�Kni�2#���"�궮�^�eH�˙Xi1��~���A�
�㼳�Z��j�U ����|[޳WD�t�s�E��lD���Ȳ/;
"���ړ?�N ��7����ۢ��`�5�y�!w��!޸�
�:.p[�K��k��*8_j!44w�rT����>錤k�HOL_ն��"ˏ��l/m���Sh���YA`(Ɩ֗wMjh"��b�dF�if���R7bb��.��YYif�B�s���*��
B���R43���K�T�v��6�UY(H��#,�E��x}yrl<s��$g��P�����N�=����&��%��u��}^�z��b�Ym������̚B�z�|1�Ғ��k`mz4��wB�baz3��sN�y�{�����p#��VZ�����yMLM�:ϮUܲ��Λ ��V6����zS�/��e����xe3f/�^fA�+R�G�����j��D��E�Z>cMD�.8��5yX4�
,���p ����Nӂ�
����?��KW��@��ho������l�{�Cs[��wङg#�T��e��N��Q��[gi�n�QeßqQj@:�|���j}�b�Bs�j�gJPu�FIS���xsy(�tp��C��B��)otf=n��ofc(���l�s?�q���p�"�?[I�:^I�la�0�X��k�gآ��G�?�^����y!ϿA�t]��G|������F1=���W�;θ��U:<P�� P�q&�%������m�X��������Nh�u��6=��_�`r<�-$wrU�����%Z���`�!p�w����j�-)x��+j\���?���YY��_|���\�GB_�,�M��h.,zJ��)T� 0��=�m �Aiz����\�X��/�V�J�/����30���2U)2�e��s׊Y�s�q�u~����^��ߗ��ZS�I����ͫM�ĺ�y��h�^޲�������u��1|L�Sp���2�AV@��R3�
ao�S|��Z,�f5�b����<9�	�6���Kp���X[#�&�^�gͯ����H��n�㍤D�lo7�X�O��U�_j��Ё�d}Uգ��2���L���D�~�O�]f3�����(�N���%�܊c���y7��>D-D`������(�V�-�NUO3T�Us�ģ�7���B��/��R��2�+'�i[d
�ֈe��@�m9@x�U����(�`������2?	(��r����g�[Ze$��n�����ë�}�a�$�Gv��뼽#�W��J�9��e�sCqM1��hz�X�ߢ�=F\$~���e�ئT��ئ��K�j�6��ӠR�����a1��hKǷw�G�CF������~K�0�{��zE"$�4U�	`�����I�zŜVt�|����nOLҙ��5��#�$*�ǵ�0��sk��r�YN����"�3_���SP��#ٌ ���,��୙�jj��HW���:䳉ɶ[- ]�i>�6��*�U샳f=�ِ�Է��U㩈;T?��Xr�ڃ�a�7e���먝�X���Z¯�*؇d~�7�7��,I��u+��4�$�]%�A�;���[�f��q˙��%������F��6	�	Ħ](����k�[�Wq|ʼ�S䊤����'�\Z#��Q���`���v�,���R��3}�,�Ԯ��=~��B���6��I.��Zj���eߚQ���?��@�[<���N�S}�=��z���w$�/�H���P���%�(ꥃ6�ImK���عPj/Y��o���#I����-"]-ꇋ��㌳������xLD��ܑ���E�n�D��V�>��9--�wF�X"�fw)��4�w�K}}M�\%�eTNn�"u��n'���o��w�XC���>t�����s3�(�����1Y5[�������_����\˗���f^i�uSw�%�ʓ�Im���Y���s$��2��Vs����_gg(22]u�/�>�kY&K��3��-%����ף|?0��pqG���r��Ɵ����"b.����u�>�bV�h�P6���zCU'�`���i�vT[c?]L�K�_X�������������ಲ��(��:�z���Ĉ�D��f�g7�4s�0Q�FzA��B��fW�f��w;�Fv��� hq�A.�T�L=ϢWQ�.W�}%ƴ.f d/i�3�ʙ�&��l�YZ��%(� �ol'�FI�\e�`��޾,<%�&v�75AK�K���A+��0�j�����J���;6�Ť+w�zH:,�F~N?R�x˗^N��pV<m�/���Pw�;:.��.��i����q�y���bd<O�n���G+WoV�5�<��>vE�դjo�޼b!��˾7�d�Ke���4P��  r:��}Roδ͞q���W�]�he�PtE�>���G�ʎ�L�*r<�J�Pe�~�_��L�m�h�`b̧��Y�~�C/�N���|�k�Y�Q��cB��F�����P�~�Y���	�kd/��s;�j��;��d
.�96q7##6ǣ�<yY7q��}�r�=�J&hF��L~|�����9G�$�Ej*@��EK��!īySK����3���W����-�4k+/`"�|�Q\�JG�9ZhlX٢>n�P	ZP=�RY�>J��Q3t�8�4��;�2rWv��V�平�_� ��{�0K�S����q{d���M��4�I\[X�<;4D,��T���{��AH	�!Ϭ�#��ߗ4P9�!��y�4 ��qUe�f[ǎ�y�H��%.NXV���w�ޜ���;�-�z�kr�k���ӄ�k��I���i&�|t��0UHe�iX�;�:S���O��*�(��]��Np�n'��u1o����h�0W�e�j��J�b�<N>�V�*��.Y^+�U��6��1.~؝E���������q	ͷ�.� �3Μ.�ϱ&V������̓�<�bE_��t�n��5��?��"��a�$��X&���p�����fM?>
>���A�3y������jX�W桉���+]6���] �{J��-@
ճ�==�Z�;;�ݟP�D��Ҹs�������|���r��lSfɵ`!�b�0�6�	#����R��_�����p:3�"��W��S�J�~�s�ISٲ�_���7]�cI�b�b�GO,o^X���)�A�W�G&��bD�9~�8V�v �$$R���L-�8�+��,��*3֋&�\Ƌ�Gw>�ިH��ӧ���h�K3�5j5��9��;��p��"����ͳ=r��gN�1mU�'Y���m(��D��ꩱ�GG�Cٕ/l���vUz~��_S����G��X��Ҿn���:-,G��1'p��4�7�݈`.5`�"���6���0�pE��u��V�����
���q��-ؚ�;��uA�K%*v�Z��"ws>gS�P�%��G�V�6��Q䅗�`՝w0�KB�o�t���HN���9F��O���/�H�F�����Cᖄ���,��̹�W��.��O�aW�J�`A�a݂!I5�*	)�XqxʾK�?Y����?0rH�/IU�=�}��O�@��Ly޲a��~�w�~�F����]�,��|GU5��$��A%�{����v)���ʽ�+�����2?�#>%sO0	Z8/�A�7��`�N
K�^� �o���i�Β�QX���ɲ��+�9����U�_�4hB8�t�`5P��9n�m�5��������H	jxu���H�6Ȼ�K�����]I(C�a��A�o��e>!`f�����k�~�SU�tĖ��3]�6�!�}�Yp\�|��ž��g\�n�F�6��ۺ9���ʚ��ȡ��_nEs�S &�%)���Y�zF���e��o3��d�I�����J��5t�,=�q\ ��߶)�WBB�ӗ��;̵�o`�_|�{h܅{R��6:齩y5��<�3{j�[5`ie��԰��+c��i�%�$�͛���1N�*�oywd��&�X�)�tH14f�E��C���4H����P�Թ��+Ū|���(��`��=+F?�e`7�[þa�`����.�gA�M���QY�[yڭ9��u�����gQ4ހ�S?� ǣ�8e�Y$�{˧�f.��9�ݮ���Q�@��~�򟞊�?����vn����cƭ]y��ROQ�VӢG�ߣh��2�8��f�w?�Q[��c/j�P�\�"�B���>�	�x�e'0�캈\�U�^:���-3xζ�3A=��/��a8�>Hv�c\$��-ڗ��GB`?<��G���s��=�E�y'�&%j��]��5��EW��}0���[�5(������]!|>nBq�Z0�W8����MM���yg�6Cr�6����eI��
�9Z���
T���o����xp�����!�{Ofd-�bG��$gj+l���j�ޓT����'�6�s	���� /DGަ�7�u.�{К�-:�{i��{��fV��<������h��n�Y�3�OU0�s�y�I���`a���NJJ��,^|��b��_Y�b���.K_Z8v=��'�vM����� D�� M_�m�_ř��Bn����+�{~nI�SMd��1�8�L��d���QL���Ԯ9X��֕���E��'%䘄e��Ec�	Ӊm��/����Z8�5�0��F��'�Z��W*���?����b����F��b���!����e߻]�ѵ7�41>��t�A���Q]��� �%	��3�����k�������M}"t����~[�����[��؟�x1q![ݠ����g��_��+Vs��N�$l��6�W�E��ٮd��t����_7�,c0J��I�+��	�K�W�5��wK_�H�
\?]��N���h���/R��� A��m�)lㅱ-��.6�SbT��N+�fr(�@�ғ_���a�AMQo���
�w\K�cF�~�k#�;;�����[_H���n��H�)|_/bS����A�
�EOrX#�#��WþM��B)+�ۏ���`��J4�1d�[�����iR���P@��d��I{?9�#Fm�nM�>�� �X�&�h�G��^�g�Qf6r�)8`ER����fdUU��Ԑ�����W��8f�9��#�(Y~���a���_���Ic�X�/T}��$rKO�c�Iv�G��s��1_>7?~�g����D_�
Se�2~8MWI���T�p^�z�s�R�d�>�?�ZN���rߴ�{���\o��i{��	��^�?���z�"(+Gb�N��0�v����n�k���2 ���C0�迷��SZ��I��|
�]drO?�2���M���e�:��jH��.���v:"c�B@��:�X��k�~Ֆ'�ݢ�o��Q�������)�^�J�ק�����L�0���~cZ 3n�A0f��4��iiN������H�H��d$N_qq�����C{�1���=O�:l�<^g�@�pC^Ɔ�r��N��J���ap�œ�R��"�w�����Pxx\�r���}�_��>r=zm|W�du��? -�~�@3�2ί�?�Y�"��7gﱱ=Й�%1=������?��i���?;}��l�O������߈]���aY�uce@��C���� �hz[���f��{��g�!x��BD���D�$>�z������C��(.�v��O����I7�����(sa|�)���l�u�!�>2��Ά�j
@E�tZ[��Î��}������.��DQ���a���;;�
-9��8R7���O|�X*��Pk�e�|▉��x@��UO{�qCx���(��>���!a]�?������.ɐ	�c�v\�_3�O�+_
�AZ�q�G]�&�.�}�D�d�и��"����Қ�ޖ���GxĈ�#��q9���2���eqK�h��3��L�.g\��ۛ�Dź+@"�˼����i�b�e..�,t暹ήf�Dޛ�k�׶����[T��BWk�}�$��Z�����}bcCV��79b]���!yg]z�B�惑�&��*&����D�f��G�-ʥ���ްkӹ�ا`��ءWs��QOq/6�K�Cu3c�$����1�JeN�jp-�(w��vj��eV��R�vJ���	��b�J�lH������/-7M�c/wl`�
�.��ԽL\vL83�n(�l!u�����{|�3��v�Ð������q~��nh�_��i����߼7_���.n��P�&%���;�)�_���R ܮ�hM�ަk��4D�����<�f.R���,��Y��_v;�u[�XN��L�j-�)�f�a�&�y�'oV͏j��y�����A�u����~�#� ў��[�l��"�2�LF���n8��!6b��U:߆5zCNC��Ku�A*'�8�w��~�2ϖ���{��Xp�v�Ӈ9t�<�Q��橭芑Fz����я|�;ײ	QAس�K��+/�3�,b��*T(�p������%�QI��$ ����#k����l'لݏ�U��"�NW�Z�x�J�X��a"��nlq�y�/`�޸��߰)�!6^,�O����zQ�6k��K�KV��#�y�}N��u�R���|y`�{��O��;TC��������5� lWr
��LWT���Z��u���%I�Tv"��D��`�?�gt/�q~���ކ�7�u�]'��t�g��L�otyf剌�,�2z�<Q����9�2�ϢҬ���`����j*4(�d''��ݱ��d#�ȢX�y�q����Th)��+l�/x�6��^D)͘�+1T�o� ���p��C��R��T�]A�b���6gI3�ӯ5D����n\�4lD���m�+"cU0up3N���?�����Y�������W�{���f^w��Dǌ�ޭW$�02c�M���mm%xR�W�Y�0
e�<��y����7���j�KZ���e�-�ӥ�o^H�X�Q�BF�]�fM͐s28)�)
��T���RA�TGe1�.f��hkĽ9ա�����Hnġd������$P���m�\~��)��Z���
��W+9T������������tf�>�����m᎗�i�]�qa�2W��Q��d����V-���f��(�wKo�\��	�T��'���R�D�b��6T�<mWc�{q���QZ�P� � �ӽ35Zp�����-�5����?W�	�>��� Y�*�63P##���c�dv�����B��B�@s:��_�yy�� ����V�ְ� �WH�Hs�����_N|4c�t��A��٧&�7��m��@�d�Cnİ��{��� ��e[V��C�]/.�}yuDy��H���c9�G�,�B]y��G�����ń�/�d�t���"F���޺1�:l���m�=|���@���s��b3�v��E��+[���h�2��W��d�=�՗M��ʢ��1���^��QSXK���8���!���q���P��]�S������O{��Ӓ�]ñ[��3�0�y��w�u�b���bVLj�����ޭA� ��kۤ!L=���r���P���W����=\rk���A?"W�0�H��,.W���y���Y6�4'�����:ſM�Y�W
�^�Ň�K���;	=�V}�%̄�Vo��3q6��@�2Ï��V��i�b!6�����U�#�ڲ��M����ӥ�A�,�9(���MЎ��jb�>�0�ُ�w��:��K~�&	��
�_Mk/PLbS�����|��$��n;��<c~� y~������6������A���*�oZ��S��zSB��e����^�(���KM���R3-aE"�O^ٿ���Гdt��}c��a`���pV
�:^I������6��eW�����b�F��N�Etb�yB�%�U~�p�Ыsu`�tp�:���t����2���_�S[�\��y��T������/�3:HK��#N��$���Y�L�;�s^C�9��|[�eʙGH��N�DS~n�qE����Қ�,�K�ԯ��4Y�{B�|G�ŽeiL����#�ճX��{&	���U���1��<���1�
��N���-߲:mLVJ"���
�f��?�1Rk��Q�6�mݭ�ZK�$���KI��%\�4�<T���nȜ;�&~#�}e�${9Ǎb�7� �&�P㏌L�'�EkX�l;��u���rR+��\�˫~8VЅ/�d86Äu�5�-��#�e�1��� �A�Za�;��<e����o=�H�n��ʎacz�����ѫ�c�G4I�2{�ZQ��⊡��y�hvXIQ��w���C1�J
i@�wVa��ȳ��M�|?�H#�@��c��t\�r܇��z���鰵G$�-��=p�v�~]a�!w~��|>�$��!�,���|��AC���䤼��U��O��r������� ��7�l���v$y�_v|�^�EW��6�G�к�r�4�׌���� {��Z�_�a-M렞>��1�������L��^ڕ4����-Ԕ���z�@H���Oҷ�b]�+�ǳC�F��H�᭱K�/�^Д%�!��Fj[���?�A��~��g�p�<�Ƨ֣4nFY�?�?kd�x���\߹>G���ߢ+�=E������r����hyO����*��Ö"�_(�l��0��(jc�l����]~�H[%W����	�`d����&�R�l�#�W��P��;�`j�i2�v���ޗѿf�.���7Ҍ�9}4�{�s����:4򭜑a.�e-GBW �W�L6��ڑ?3�4�^�>�]�i�2PA��E/>��ŏ�e���{E���� �=Ğ���m���ɧ����W�1�5�� W��o�E� �����h��t��D��o�*�rh=���眽U47���b���q����+��Ȝ���lq�y!3�C�{R���j!آo��	�sp�9�qx��������UUޓ薾[8��t��K!ޱB)+���p�d�/�p���Av�~\�϶�*ྦྷ�u~�;2��h ^O�	��jo��!�l��tlٽ/�]ri���$�fߺ%�F|�����/���܄��8O�ZfP��-Xr��v��~�;WQ��Q�N�.]�L�'5�桲�ͽ�M~fi���5V�F3�;e��i�����^���Wz��1Q�-��?r��u�S@�p��Q4[XBeS�t=�>�?\i�&g(P��J��E*��s�)I�e��~���*}TNM9h�Xo^����僲�jd���	�a�F�pH�K<�g�u��4ƨ�M~m�q v�3��k0�\nEC w=��ϓh���g�H��"����3�\�<�R��js��q����:=������q\g'���;��|[���n�}O
nC|/QW����9��ZJM�P�i{�@��{�lt%���b�l}�e���)�`��{�U`��O"20�m2�i����l�Pj��f�[����J[����Q��K��7�-�e���`DY��?!���R�s���7��鼖��������Nq�G��f���)�6�Ṩ5E�}�J���f�y�\��J6n���J�ٟw�T�+!Ӕt�����sjV�`A��q4�$f}<�mdG�K8iOb&���֠DR��k���O'
n�x/��ss2�xCS��_�:,�H�!!2�_��x���/�t�_�*��%tu��J�����x"����R�"FH�F�`��k3?ai�eU�݊������g %PI�$��*c��u��fP��4���Bp�7����ܱ�r�����sV����+�Qk��}��I����� ����)�1H#�Q�����ӓ�&q �ޔ�#�s �ČAڡt;K|[�ʩ��Y���g��n�T�n�è���w�Q~��#C����ut{��<j(
Iո�)|)ۀ�gT��4��!e[�������Y����G'����v���Ϗ���y!�N����'x��H�|ܜ�i�H�ٲ�M�kM̕�2u�.�p��?��W@-U3��r~	��W�Y6A������1s�	C������_J�l�֭����[�i��������*�1����$s��}hY@�1J�<�ЦɎ*��1e�}2L�>&��e�c;�nz����e�D^�p�"��ʰ�$q�_wk����"HQ�*���(r)~���$ϧ4��	�A�9Ze@�����z-��Ԏ�NI䡣8���B�������G�VC�3�=_��=��:��`� 9�N_�����0&Ԙ9cz�x�l��3xwy7���ꌃ�l]V��t�j�����,�qMX`a�/�?�)<�x��x���S��w/T�6���S̈́`���{ ǹ��y6VL<aL���}�a��-��:���G���۾�tl�E���8�;۝�~��P?���Y�C�0�U;Ÿ3��L�=Cx���s�s�&^�
��͹�����v@ٮ��;Y.��	��Oy���l�0.���\�\D?-s��`��jc�H��@M+j��;��V����Q&t$vq>�k&6Ƹ>GR��P1��o��h��g).ƨ��w�Cl�oǹx�3v%��sNɑH}����W;����[�����j
.�)�m^�HL���a����(TN�lMh�춹9�,�i��6�I޻/�%Z��2N˒���}��`�mx"��!���"�fƿ�n����AцZg��fC�h&h�H�)��[�S䂯U����g5�� �ij���zsx2��pv�]��o%"2�"��G|��WGvuS"<��u`&��U?�BG� �^���o��88��ts��X�9cj�C�xm�Im��3:�Yns��Z؀VZӾW6�7�
�k�̗�Yڄ�J��K`^��'�Ѿ�������;Q$}�AF�W(��1T��S�Q�@w�,��P�*/-S��|^��)\�J�?0̪�c��ܳڿ1��c5��;f�X�@Sڏ */\�����q��OU�;Pꐼ����o��Ph��1����@M$X�
ʦ�+b8d�S���Fg�S�\�}"���#�b���זk]����跶���V��dx�Eޚ�Io�پ|@+�\2�r��������be�ܖ�e�����^L���4�^]�C��-'�}���[�=g`�j�[��!n^d�u�\�4��=V2�4�lI�U:�;����Ѿ]��k��Pe�G\�Fm]�*��j�S�ڻ�#-��y�o;����� ��u9}���|�r�K�Zo�O��e)��5���R�?�<�������b��`< �<��˙��c�*u�ٔ�-ݍa�c����b�5o�4~ס	/���v$N864�t3\tv��t��U��+I�-�C�y��)J�|���vA��� �}:�{qg�[�����J��G�L�U�Շ2\��Z1�ͭ���ȑ���u�ʃ��mi۪�d�흡�l~�ي�΄3����VSZ�OZ��r�e��W6Ƭ��ϔO�!GŸ������:��r}�o�z5Ѱ;�ҫʶT-�q�á�3w����x[&Si�z�/8�Jx���PZ�s��r�4�yz�Usc�;f�yܻ+dj����^��������D"�9���y����ǅ��.E�ї���Y<��9�k꧑k���o�z���:�{*깩̙���䛶&J���G��I$�$�)����Ez��jr�t��,<������8	wՇ	���h�߇ن6W��ѯ�=�ކF*������v-������fM���|s,�ɺ���K�8�H,b�"0�ڪ���lJ��R\3�>s���箒 /DKO���r�y�{�^�mㇶ�Z��/�2�����!�Gڭ��ǁ��{,:A}�R5%o�Bk�]=|?Iϔ-t�-�,�ꏊ��칭j�x,Q�F4�{����c��S�DsXvw�vX�Z���o�J+A$C$����8�w��D3e�H�A���������i����'~*E=���Ì`�%����6v �'=
%�gK�������Q�}�Wԓ`��_"�5`�Lǯ�n]�S��Қ�;~�h���1.�:R<�펼��9>m�im�r�ɕ@��&��k~���&���ի 8�R��+��w�V�=�yH�F9��"�S*��)����i�[�a����A������+���iuo(�X�-�C�>ĄnINF73#���)��n^�LD�v{��c��[��0F(f,p��b���ܫ��؀� �n�O`7IG�Ѧ�q���ᤨ"�V(�\�Ò���I=o�ߘ�����Y$N��~�*�O5�`��]�LXn�����R��h�q6�2?T�xw3��#��j�ܣ1@",]鴓�
�Ǵv��;��E-�y�M�˵��u5�7u+/�v����J]ld�u�"�`�B�*��^����1qO௩"��$�x�M��j)�0�sB�Y6>}'ΑY�.��7��[�q��X`�l�
9MH|�t��f�+��>�V�$�Xo�u��l�v_1�(��ˁ��}[`�o8�0-}�k	axG��Ƨ����x�V�[:��C�E�UFj��Q�NsF�b���Z��x�MN�ĽV�ݥ�9\%rJ�p�r���C�w8,9�����N�w��|�h�d4��4�����e�9�Vw*�9��uwW�=H��E�J���j���@B.�'����s����2Q��bh����ũ	�z�فҁ�S�&�K���t��9X���!��1u�s�b_p��o����C����誢�X4�˥E��o��;0������Nǅ'��:�KO��;��U��dUȱ���`� ��؍���i(I�Ɨ�/Q&�և��nd{��wqQD��U�cy�M��{�ߍ8N?�'�v��g�������B�DY4З�?�J�(�>(�T�ͰI�u�0�s%E�V)�S�⸌��������1�az�� ��r`�<ʙ7���}K^���ek		��nZ���W4+t.cH�C_/S��[�u��X��$���u%�yp�h�0��O1��s�m��K-aȤZW��F�4Q�%��!��*'4��e�Tv���a�<�|6����>~�9LwS��Ǿm"^I���ҵ���!�y�Sy��J5m=��61�ħ�D:a��z6%+�cl��7}?�q����.�~����/⸛\��mt������@�E*w�T�+ �����h7��lJU�V0��8(����~����{m����9�S��?-����|TM��������V����Wb�]�lk\��7��5�9�2���έ�v��k1�7����J�
��}MU�r��#`���ǽ�����[�����#���7n���s~�#����O�_}��Y�KQÊ���#��_l�׷�	�����w�����n����U��\ܕ��c�/�Җ�A�ɏam{	�P�*��}�`j�f;��fC����A��}A�R3H�����l��;??��������
�+Xe�m���O!e\ �F4��`1�d�obސ���f�ٱ��\����*T���q�0{Fؼ{�<9X�U��e98^;	ѥ�#�!J7ͣ'pi�#�n �/�Rw�FJ�{y�ܾ�4eZ��st�ibX�ɺ�bs?"ל9�\s�!&{`����G�_>y;`:TG`?P��s�����^V&(��n8I�ä�x��U�U>c�%��贯�-f��ط��)u��/��<i�����?R�+�*9�-��ߖ��N�\�r��B�Z��I��ABF<)w̞"��*���_ל��h�R��t��ÙR�̳å��Oo<^�;204|����50R��V�E��/G���tڵ� ���������-����ϳ�~b��٭+"����z��70��Y�%�}a��ӥ��{*F����x:Y����e{�հ���Yon�(U��L�Ur�!�$���Ӽ�����ք):*�;��ߡ�+��%��T����}ض3ʾI���	ޭ�������͜Iz*.���l��FJG&�V���b���gH#��k���S�H����uy�p�b�,~'q���.�*�N����M���ax��t�~Y�X��筯a.-.��8�I���B�re���ale�y�&H	����%*#���oY�?J���)}���+�>U���)��{y�~c˚JWt�_�헺+@����8�4��50Y	���U&�9�A�s0�,���퇑�s:�]�'ŭ�����F�X��}���L97*�m�ٞ�\C"������s�������b̆�͘!j$z<�r������t���f���,|�e/Cv�vP*o��¦� f��jM�_�_��P���V��*�7�m����đ�����9J莮��s86�������/�T������-��ĳ�#F��*p�zD����em5@����-�ęJ��>�*��żNz�d���}���N�d����h?����� }�ޕ���%��=FP7\ [*�\���#5m��Uې��PW�`ˀ�Lce���	���H*�c�-��_�>�.h�̺�'҃H������A��~{�|-����a�MǴًHg���	ñ��V�Rp6�Fm�?4�WP
����(�" �c�
(=XA��H�DD@��$�J�A��T@D���B���C/		%��B%�{g��>����?��[g��4���d--�7��x!��M[e��ع�t��o$�/A�J<�]'�t`w�/C򌍟��n0_�6��Lnw��w�W��5�)��3՟	\�D� :� �V�+�.�C�A�$f�V���\Zm�'N=T�F�L����ՠf�\	 M�3�����:
W�
�̓J����[��Uy�Q
qǚ�^iA����y��0�VX��]��Dr-�+��_�j��ݝASW	q�������-z��?؉��J�C�K�}��,k�O>�%����9I�1�Dt��rbV���'��'%�/��i:V8%��_�tj���y+D�f����Wb���knO�*��Q`�?u��&�)�̔A�xF� d5���b�]��8\U$//�X;��k�E�0���!<��r?��5'���W����S�$��֧��L�
��/c^��N���k��j���DṾKI�|#�zK�����l��γ�[}V.�h$�p�n2ncT�^+�Ul��G�6st�8ML{� ��p��H�ٴ��a��|�	91>�D�{�z�B�#q��CE��F�V�֚ ���vO�,87��$����?�3ǫPڃ�����o�Q6��#�F��tGaȢzp��_�����z-��/ݖB��\F���p%��1��tZͬڈ8��!}y�9�[����muBJf#��͊dQe�%���u���pci����"W�]*s�\��iF�*5@ۮ�X�4T���Y�xJ@W��>v���Y�������A���}Khv�x6�k�`�^�Q�^nً�!(7��k9zz��nфP��zp6�sp����7��Vsx�v󉤒�H���@�}9��0�K�՗z��e���
��X��i���%�Q�'lEĥ��-`����}��$����ŏT7��H�]a�K�z�v���-LC��@���O,5)�{/&�Uձ�*r��/�Vq{��#-�����_��3\+t�\#���ƙi9F�LJ��+~=eGZ5:tڜc��tG���w�Qˇ���mSj��{nx���N����a����E�:tDkʝ��ہ
���p���`�����ַ��)�}q�Usc���cf{�f��QF3�/�9��߻�A��~s�3��4�����g�R����[¿�d��C�Z4��7i)�oM4j�1��������C]=f,�e��`��
oe�E��?��^�m*��(|���0Ȥ�6+��JQ
�ڳ�<�y��3�Ɍ��_��)]�Ou?o�%���Wh�5|jǆr]�<�&�|#�
ƇsTis�r�3�}Iȣy�� ��p�'M��Ř�v��������c�|��{q�s�SI�N�$O��K*�@U��d���K��&��hAꍳ�m�}���nm�e){1�f����z���G�[��f�#:��f�>h�b5�%�N���NE��[���?U[��,�4��{�ׇ�=ӹG~��Пt��~�-�2�u�[��V���5R���E������y�Nk�J�����Xn��C�>�]����k#�HM�ێ��P�
���$���-I��>c�Y#�ūFK��������yi�O�sהw&3\�������wۭ>Y����������Y��⒏�I-�����ɮ�R��}��o�P��	o����Wsy�Q���yRl'���+��}���܈"�\X"�t%�7��(��!�9W�ȇ^�O��z�Tl��(��/E� �LY'��h�$P�U!��%�[RW��p7$Y柊��:O�<hL?Yz�Akx�.�+;b⼐����>���q1���b���4+�I�M�ȩ�t
��Bhc�א����ʷOʖ��b s*3\Y&%�)�)���-�����5k��,^g@��� V��	%c�:�k���<a>�/ל�;{|�'�碑;ll�4[Z�L�ld�7�/�:��,C3e�p�a����P灨���vJp����HX@y+��z�N�5i(��������.�^�?9����}���Cx��:���K�{��$c眏U�:��+�_h��s���?#8���]X�aRc�Ս�����y�Y�%rX,���kD;7@8��'�vV.PG$���������G
�����1�F��a�b	d9o�q�b4���n�a�����e��{�['��	�@)�ENߐ+��VWzy��ϯj��}�������3�V캪3ayϿ�(���
�({z~݉�D_��T�^Ih\Y␣@,��F��h���И��6��ӷ�F�Q_�C��C;lo�鵶��|4��|�8�X�1皍O�5c�-�����M��l	TH��}�!5�;�s!�
ZX13�'
PN�A՟$����Q�R���-�BX>��ͦ�_5Ix���sh|���C�o�ζ�ǎ3C&,^v���_O�ÖϋڅD�\�x64���ɶ��5����^;F�u02-6��!��p��S��`-�f�ܥ�Ⱥ�y��O�W��GLn����y�1~SI��+NC&xߪu���>#-�	0�nx!�4d�keÙ�.���Nɮhu�����S$_ �^&$��a�� �c�7�}����g=��c!�m^o����E>hj��2;��F9������/�V!<�8�����:0��9&]�)|��o�[O����aR�o)�{L$z�:_-�A1y=�F�ͣn/��Մk[M?�WH�Gy��}�ӒNJ0u�U29���|v��7�����  �k�-+�W�q����~+��;v�,��ъ����Cf*��Z@;���m�H����Y�W�mU�5�x�=������s�V/:��ϛSfX{���}���'f�zNQ���-)"q�y��v9D��A��s#d���N���E��C��`���"t������G�U.ޒ�3��~�`p�(J�7�J�I�I����=VPf�S���T�����<ض�����W*N��4��a�"}8<��gf���Q�:h
�⣯�T�sJ/o� �],/��n�붴�ݣ�e�(��_;��hM���"& �)�*ʥU�'M�c�ü)i!uG���Z��0�t�9�M���Z�j"F���<!dh6�`�O��+���}8:�9�����~����� s��x�yg�u��_�#��zc�[��c*�s�|��*�p���Y;��0���� o�i=Sm�_2J�%"�s���^�|`y ��D͹� �¼O����5�
\���q�����m�t���n+��k}WX��X��+�.�	���Ac%�����3wY�g;�[�P_��{=�{^�9�{�3���W��S�w�Tb���n�s6d�$������\�������/����5�&�3����2�i[+M]%F�G�X��/����S��PE�N��@
��uU��fS�La)KYg7�.'��^��v�M��B�x�u0��)�k��`�I��CKv(�Vk�r��L�F*O.ûh��n(i�RRL:Z��#k_vK�t^1A��<�W�H���ZH_WIP	�9��=	fa~G+[�g�E xFO�0�m�7~�u밀������+ٰ�Kq��n�w�ͭ����|��������+�HW������n��P�^��}�w.�ư�-�s�k��1�03��r��pV|����������}I@���%gGz֫���=���D|$.�����}�7D�	<�/L���E]&��ѹB^����[]"I6��a�G��j�^ra��~�V�G��U炚����N��?J-�c[��{e �)0������_ElS甼^j؇���j�D�.݊9�"{��!TZ��/E|Q�dR*��0�X��t�\��MQu���r@9���~�D`~H���*��	5~vW.^Y1sw;kI��5����r�����>2������ 2�?���a?d.ȣ�d����r�`��k0�#4���1�RV(cm#6*ʎs3���5��Q���f�{x�L���b��y?fBf����������P8� �posT�v����5
Z;l{�B�k�V�F�f� Oc�PyH��p���|v�]o5h!�����7��M�ߓ!�B���/�r��UU���ߨJ�z��i��3��*tzc������E�5�������)��Zn����<3���=�:������DX5��]��;34r`�'�t�W�0~��ԭegl����~B�����\|*mWa��~&	�ă������q��^����BӁ�y�}�M5�U2Ać6E�e�M5	z����b�r���&�H�A'�v}kU�le��4��J_h|q����`����}�I]YTb��T#����w�!��2�.#�� �Ӵi�ÕͧƓ9 �Pqt�ԂC��-��.[��H��o�N��1�����y;3f_L��7`�]��A����X
M���+=L�����Ի�to�4LO�L~� _�ͱ��C�z����؀����<�:���t�x����y�})�t�d'������՝�!��QҰ�Or�˖#I1��q	
"u��;��(�G,��\��Rť�@'�]���v�s�p�d�I�}�hYe��-8ue���<z�R��� s=C�����o�l�`PO;���[=@��P��9e���'W�iQ��O̠���Z��U>K��O�u��Z����`���8�Ŋ�	��z������~�۽u�7ox�q$�vD����k�{KB�_�Cy)����i L�m]~؆��
�K�.8WT���$[�V�K@�Ս��A/���K�����zu,Nwa݋e�i�r�c�o5��/V�6A�L=��"�Y�V�����oK�3���1=��U0��T�*��db����*�^�8޴�Z{�@�f<|Թ���^�u�A�"��U�9�iH��]�"п�@\T�N��ՐWfR��*�[�b~C�R�����G���������au�:i@�0k���� ]�#0�L>ݷ0C=7q��P'mY�����U.��*	i�u8Q�\X�^ĹMW���H}�}�~��I�T{.��;��\�����x��a?y�8�ަ��gum�[S-����KY�dK�r�iV&�K4Rׯnߜ�~���Xڵz�I�$��cp��_���4t��V�8��wC�3>9�b�0�D����+Џe�y�Ou	�$o�-襰��5C��Q�}m��TROd0L�\V��/�T�JcA���I<�A��VRѯ����H�H|EH����8���V��X}M}���EUE5NB�:`_��$`��N!ʒw���E������UV���qJC�����]�o!���3vL	��r��ڥ�I4���Ϲ�����T�'r�U����v��3�akKE= �ƛ )�k#Kj/�1�`u��L�i��}+:���T�uF�!��Z�1[�
�<�V�=X��$C	���ݻ@�^���� %�)�3YZ�
 �A�bfW,Q�ٱd�s���
nS�b�iX�f�"������>['�����׈��9Z�0M��o� �M�rT�f��&�~碩*
����{5�i�+	��g���m��a2���%�'L������'UO�y/m^B;'����p$7�����{�b� ��A2�0��K����4K�V7��QE!��<w/y��9��Q1a�f�6(�5i������-�m���FZ�1��q�:�aQeL��P��6��0�$���
g�qj� :���'H��������>�++,Ӻ�4ŋ5	Ͼ�^��R� jU�6#bTO?�>
�
�|�h��}�hdۄ���y���(�b �D����hF��%�eDy�b���9P���@-_��)�#+���sa����G��s�~t��GdmX�C=�n�{>-�5Q�j��{�(��q�B�B��u�ʅ�x�m�,�kk�eaG�+�~���0�".Ƥ�;[����.�
�(6��C!]nW�+K��i'D�T�9{�
X��<2m�*ϫa��������N8���j௤jV����c�+}����h�%����)'J�.Di��M�9,�t��Ŗ+�;�Qg�w��C�9�z�lV��=� ��:���+cw���m�	NS��GW�J�?H,1�1�5a�TU~�� w�R������ڬߪҸt�|��C�Us�zp��E�2���`�.�%���`Uӿ�e`�p3}xZ4�شj�''�|�X�P��g���!I4� u�~ш9$OR�a(a�����-5�����[�a��6�Z�BBS�@�|3�����cms-R��⤞}�,�	�,}ؼ�/g�L�cݖn*j#5׬�u`����K�J;���9�n�a��pl;�xh�"�H{kO��3�l��n�D�c^b���˞p1�����)����V\9�Ҭ��U�P8�}/F���o��4����ѡ҃h~�����x���F�	����s��T"���&�y=,�mWGOv�f��N��݂@S��h3�?��w$���{�Jt�9��m��y�ֿk����vq�.A�*���9\Y�J{yB�4�L;�c�������W�B[b 	��K%����ۻ54�A�YLAE�	&��"���: ٧o�{}�����>p]��u��=H�0V���9
��Fd�M���MT���6{`΅��ʚ�ƧC�=�֫�cl��r����r�]�q`P�1�t�S�sp�A�-� ^��a\%>����-R�v��V�i]�k��	d�n�ױ���!��X'�|^	�W�x:�PYg`�����%�f\�ӈS�j���.^��m s���Uԟ���6Z����E����v͇z��h� >�dm�X�QtD9�T��\�����Bk�(��a�^/�I����He��O�q��?����S��߫$t����ߖj�����^���Q�5]��d��e����j��H����P27�o4T1��-B@{��thZ�9a��C���U�{��O�����o_���%�����Q��e��h��mh�����)�S@̀P��j�ݎvS��9�~�P�x��H.��iUCf���9��~l��r�\�N�Q$
%[���a�!��� ܇ P9�}?�7�Y��ۘ������5��,Ȟ<3���f�d��:��4}+a/W�#�d{�ᎎ�����8&Uv���X����@@+�[F9�:�b�������k�RW�]�ϫۣu���O��m�C��gf~�_�@����`x��Mb��J�hcᮼ�"��]�n�z���]�ԝ-$=н���wo�X�B�� ��GN-�H5��<D%��SH�|��a��<ˤXV,�޶�\=�ۛ���,pX�[�w��iF<�|�����}�u����(݌������9#QGb��$�겄-�k�R�f����D�i�j��*@a�C�S$ل �q6>2�xzO(��l��Pg�օG�u�**���;���[�g��`,�Ѫ;���l'�:�9��pv쥱s�T(69����q�8(+����6�%GP����W�|�Z���d��V�]�]���k�� ���f�pҖy�����^^.g����fᥐ��.�Ǧ�-��U/°�̪g��a���:!I=me諡ަ�M���"�L�y��g������`�O�헏0�<f}�`�}���fJ�e�c����n��>)l[NF�E�������2a!�m��u�;���$���҂���D�6o���p�d�	0����1����1ٹ�:�������THقu*�L���^��k��8\�͐�$�@)�ga�ηzɂ�7�;Ɍ0Sm�x�ل�e��[�L�c�d��gݯy��6HKfT���^��*��}D�$����ʇշ#Q�s��E?	�j"V�ޜ�־��zf��%p����W��i_عV��(�%�*P��}����ט�sG�W���"ʇÈ:���Ie��\�n����Ƚ^%�)>����k���PK�6/|��RJP�u5��%�k,� �^�'G�8R��f�dM7�X� Jl����Dxҵ�fF�0�*g?d
���i.$�i�V�&|�&� io���\�w��hE�G�[g&����=��c_�a�{�D��o�=�I���?��ń�t@��.:���7PP*��j��B�P��9<�<���G�,��w\�ɼ*|xe���x�BȢ�]+wv����$����K�#.�mdM:�n	�GIa�b2��?�K�)�Sz���ǔ��S� ��epꤷR}JZ���M�`ʛ�hIH58
e��]����J�_.<���{�$��1+����TNm[�0hZ7��w0a��#��w��&љ[�y�CT'�J_f���zZl��������Ra�VE��B8�U�S�f���5L�DJ���<t�Z��܏O��EzZe=!~��l Z|���ڻbo
��vu֪?��c6}Y`ס�Ϊ����@��7R�O6��`ϲ��`��di����P*��uU\��@�^(�q�kY�P�<ʓG�k��T��,��v�0_<-W�V�=EB=K����,�ˤ�r���Վ�@�tcT:_���<�D��U��=�����W���󖱈�Ć,C�2�o���Y���qO;���HJ��~�a˶�Hn�6a�;x#:�ιI��������T�M�"�z_W0)�#�
��5%F�|�Q=d���@�7?�~���_]�
S�f\���K綮����]��q�����1`�hyiM�lÃߩb��w�@��v�l\3��-���.����:�����i�}���4�ƛ���q��ae��bH�YZp�x_��Af+������9��'�����gK����M7��3̂7�Gh � ��}�m�� ℧��	��.�`P�UI+�%����3�^�R�0�?J�&����HZ+>Z�"~і/��[�o�R6~켚|���lsJn�"E��M\gC�ty��Wha�N�	�D��5��M�mu���k��aL����0Ѵ~u��M�Mj������i���w�7z�ɍ�=����J7��C���	D��|���m�R>~���}���X!������]��X�H�3��w��Vl�_�/M&�b���͋=2��'%l*r{w�|"�޿��c��q_��6���	�<%���$�s-
%J��eJv�?㍷,�5�K38������)�G?n9�$t���I)>`�!����.P�f����?��h�:G�H�'?�x��b�gȘI'T�w�)ۻ-g��pe�20�m����h��B8��N�
c۫g�����=Ƨ}�[�Wn���3��fn�o���!	���ڌ�k���(r~�c������O#��
��=4�o�ZU�+瞊+��s����M��(b�#���X��a�߃S��w���o�M.Q��;��O��ӟ9����΁ ��pu��7�3����Dz�O�9M�\�6��wg�Zl��]eL�\�3/F>�XpF���f��l��|a@{���z�ؘ��T�9�N+��U�=�IC98����ѡS�Y|�=�';D�����3S�sܴ<?��D�p����R<w������Q�:�o�Q�t������,@\�_��-m��T~�U��|��"�O=�|~�	�Et	DN���O�D��)O=��\!8��,F|?��X��1��aGI�,R4�C��JS"�8��4eU����
9`���/����S1��e����l�z�
���|�g�a�DOPI��8� ��5>d�p�ih�T��p��{�렡aA$vn-|�TU��笤��ݚD>�J����$?rY���b �-��4�,+qq.b|�82���<i�����ůw�S��ۻ@&�#��6�a�=�����E�ݮvx�����˩���B>�X:Q�V�}��JH���wv���..��?�%K$f|��tv2"��n����bە�&��}Qɰ�N�9�q�YY�SM�d^w���:��� �*H�_l�&43��f˷�c���v47�h�a#�s��v�R@�:�4���H�,�Ni�S ���%�3B؇��a�x�8���ө�_�K}��`=�q���	��8,�ʅ-Q�E�־�x��;Q�r.Q �ld�ܳ��J`��͙<�:����O��j~R}�z0��X�;�+H�"R<��E�pNd�3� ��L��*'��m��1K���h���F���J�>i٦��<��F;��
� �؀'���iaP��9�(MM")��儘C8�ot>m���j1���Y'�[?�!�[�M�ʅQ����5��=�ւ��/�>��=�T�-�F ��ު����xK6V9���]���·Vɶ�����Sk���?�p���Փ�_��^��*�pIb�sVf0l	�]�5�U������%ޕ��h 3V����u�.E��?:�!���	ߚ
��7�5��P}+kZ�[�9%��0��-ف��
7�:B(���b5x�2k��#�
cq;Wa���q`6�-��c��T���1>�����x��̽�����pɾ-�Y:)��8'�w޵�|����܌E��t���t�:l�2{N��~��Ar[��C�S��c����o��M�����r����j��xL�m�8�������Σa�2R=8_�����"������V@��UuM��Z�YlzHsR���\���HAf怓�3�2��0����Zڬ��NAy/���2�9.��>�p�9��9�s��<nW���"|�^��"�{\[x��uH��
��ګ���[����>7c6/�=���˱-�gx��\��B��ڧ#�Z��	v*�V�>��磐�!�?o��Hn�x[�;�.�tr�Dk�
�h�C���j,��ɓ�`y���Ϻ�������x]?�ٺ�G�!�W�?��.���Q���G>T�K��>���C��p��D��8�My��R6����؄�4Qh��x���-��/�l��.����:�Z�~x�aO�Z�X��%����]6?���IN1n��'֙�6�険t��7-��)�?J�g���(-.�����rצꡃֆ�������5F�1�$˜�����E:/n�+'��S�߻��J��B��5�/�%>hM�T��v�����S��dO�p𡚔v�Z������7��T�k�,$P\Y���It�.3]��'�;a��/w& +�&��ǙU%o�SR�p�Z��i�<�BuA��YVD�o�}�r-r{?+��w�0��]��3�~:S/�^<;����>�0�b'aW�+q����S�'���Z�����v%mw�	ȩ�Ի�t\޿:�Z��ja(��ց�
�I�ϥS��� �}�051s㆙#'��xE��Gk^3��D�/{��gD���T �����D�[m9�p$nfE��W��鷋u�-�c�if?>v=�>3�����_����� 8!���(#��t	�D�+�s�|���JM�e�ݔ��y��[�Fn+�����9���\����&oj5��o��y9���.?	��*��{�c|?4���jg�h"7�J�>w��g�ԧ?~꽺&bM�����xfr^*�`���d����{�y��};��Q�����������ť���2F�L�vwT��.���_ݫ3s-I~�5}�3��rVٲ������bӚ�� ��q!gD
���|�]R��I�	L�)��*���ϖ\@�@ߗ b������e����e��ٞ��G9�}�z���P�1���k�l�*]�� ؓxX �v��G	!�#vl�~�O���3Z��@�v���L���n*�z�F��1���AE:ߠ��9��oJ3����2<eϥ�	��ŏ��x���)M��=�/��P(�2�=h)�#���o�K�en���2�v��(���ӫ����t���Yꀏab�>����{#��~?�1l-�����Ҕae�d�]1q��2tM�v�҇h�g��9�3I�ʪ���V���RR���XV�Z�0p��Ժ��N'���vQ ԡ}qR.�q��n�\�j�$��ܻ-S�(tv�Z�	��X�,���(���y��sJ�3�,5��O�@	>�����~�|�r�����< ����0U�v����i� N=Sr"a$�`R�;�3@9g&sԶ���Lfr�N��008ďt}X��e��'9p�1��4����A�j��n���Dn��/�ɀD�8���X���B�팭�=;Zܗ��ͪmtClֈ�2���A��(u蹍��2ЍTA��O�y��RW�G�`�������T�us�۪p��2�"TMǇ����Cϟ�A�?
�4�Ҡ��?X鶀�6�Е�� �6l F�s�Q�d!N�T�o
,����z��gR9�a^�26u�)^ڌ�1��G��P���w���~ꉖ���F\WT���f�@'�귏e�ӵ--�8�+����a^(��^ES�cw�.x5��ǚ���,�j�4����r=<o	DNmoߚCQ���t=g����2x'p���Q��Zgb���zL��=fp���<�[��@W�����׼��n����%��B�%���!9��S?+��u_�:k,�)�4t�a����K�X�S�3���t��r���y�r�����[T�Y��Z�͸G�#��(S��Y\�f_x��M@w��b�.+����\Z���fpshf�3Vd�F���bw*��DCB��pf�a�U<��$�7(2�&ߜޫ{��?�,���4�ϥ����OXƖ t���@�2T&p;��金_�nN<9J�H�0���YMH�,28i�[����)1L�$����1�؀9�%��K/�}'����j�ԍO���h�M^�ZU�ike��\#�,u�Y�\�+<�z������a&�w=畵_8�Dm��ek����ͧ6�Ĩ�U������b5Qe�4ie�^=;�B���mP�f�ֹ�sf��0�]XZ���[��O7.�O1�3*�l�ȮiO3�v���]����+r�(*�E��w	r����� �Ype�fc�NM�*��4j�8�v�D~e�+v�y8<����H.���MS�~�'��p�~o[g��yC<��0}�g����#���/��h�Z��ɞ3�#��~���z��t�_�2���O8T����E,Q���0.XUh���I��x���<����J�C�NW �1v�!/u]� #�����!g���=�#�-ҧg����v��с���TbaN�QD�D�G��,�s�c��z9��B������l���[B}����#]�V?��ٔ.��V��,�
j��N�L��󊄫��kh����o���(�=�F��41o�}����â�K� ���R�7)��Y�lfZ��D {���k9��3b@�H8=<�4���'�i��(aY�`,%y����Z��q�VЪDϗ�=v�3���|gi'kM�� =��,�Oȅ!�AX��S�u~�K<��̈Ȣ)�d�޿���O����/�v�|p�ͭ����q鎍ɹmN�R�Ɗ4�xB!��Iq��8�����M����НE���-5���7�}7�Bn� ��@z���1(�:<0�]�񅤀o'yK-V����fz?�oҠ�^B�H��	���dŤd?�^4�!��������Kڔ���o�T��,�$�*7����bu�bBh}���#�q�砼���O|��Z��rh�6\�<���S�GT4�����zQ��z�������^B���u"vF�f��Ľh�Z��(8:Ld�Z���Cnz�'������@�6<S�|x��ȼ�<|�[�iG�k�i�_�����ƨ�F��������9a�g��I�����*0�ފ�Ms_�������PI�k薘P�nIUP���Ti��t�ȏ��Չ��ߘ�����8{����C�~Z���?�*Uv�f�~�~0?B��@���9�e�0X�ƾzief�����C�ķ475�A}�v�=�Q	����a|��qp��[/��8bc*�3�%Cz��}���2��#=5`a/Z]�@cc�b_O��\fLD�r��I�C����!�"�u#�7��&FN4��]���+�#���#���6��ֆQ��?^��$�|�U�Rp�F��`젿��yj�l:���9��}%�I��U���"3w�2Ȏ���l�ސݙ�%O�6�cWMk}��v��e�żv��O>�>�w�@}}�Ǥ��)�&6��і[��UI�9
df�rΌ�ށ��䋄AG��3�O�Y���N�*�^ܟ�B�|�rtL���*�L��B�p��h��+{9�s`��	[b��U}�5_����Y�&��Z8	NW">58���1{,:�G��q�� �� GGbѢ��S��Խo�\�:Z�Er�����в�Z�@5Z�!�T���M�w�k��K��۰��zJ���.�cR?ܠ-g�@8��*����1\����*�������'r�q�cD��ߐ}��z��n�F	�7hjL�v����0�����}�E�-����ת����-֥ڦ���Jo�f^�f?K�xn;y�i��-�CT�@u��r���#�����LY�����'+������Ǹ_^�)��_:U�mn"w�#�����b�1󛈮��:��N�����
FL�oS�$9� ��J�P�"o��Q���:�)����KZ���\	�mRh�xv7��HY�O)���mHQ����!	��,ɆF:&(��
� q�bD�v��*T�&{���{�#�LӢ|6o;]�NT�=���+�dA+�ݜHe}k���jH����H���)����^ۗp�$�6��Ul�O0��H��M	u���V�n�s�gB -;�<�=��.����n�d;���X���#�S�5��l���<U@/A�X�,s�u�`N}��H��G�0��.���;��*�%���b��o�[�t��1��;r����.o,S���0&�����Iҡ�.��u2\[%�5�ʄa��h���A� W��֨�g��ְ���S�`�� "��6��!��f�i.���Ӽ!�d���a]]s���W��G�`ؘYX�XoY�dX��pDO�W�1K��\N.)������n�	yL5-�U���|�������95���;�����T��C��H[F�b̒F ;L�q��fD�i|�@j��Q��p;<�Ū����ŴS� �������$<���\V�H�XCF=A�Dw[y��<�����3w����>z�M��`Sk���E�Q������i�M��?����hZ14�e�1t��y���1c�=z�d�uC��$N!O�Ռ�D��\����e�ވ6�h*��	Q��3������COW��ɜqyi/�8
撶�}�y)A����� &q��ݱv�S�3>� ̡	Y�#pa�����X�<;�g\�QI�*e��r���Q->ᑨ�	R���ϳ�"/>��rK�&���N�<�gH���sY���kncbΦq6$�?mo�
ِ)��Q�!Z�2#Q4D)�0��}����P��%��b*��������	ki	({1��`b6�כ|{n����:��'qk�8;�]4���Y4�}8�>�����<��24�@(I�ǂ��|�O�a5A.�D��~�PX<]BKn�<�]y��M�h\����\�N�UNej�B�h�U�`�Q�MH�w"�rX�6�14ۻ9���#�U�����b��i E��b<2�Sc�w�𣍀J������m�'���R�ߵ�����J=���Hp�%
!��S~j�v�-��[b��x��q޹Z��������6�{�K���ͺ��&E��k���f�U�^�D�_�]N�Q4�y���(L=w@�1����,��x���p
7&�w�=0q�h���J�wǿD�+�"3S��.!��|jJ~�ޑl��� �⤥��~���g|���$�g�/O-q�|se�{$�w�[�m�,_�=}�y���0jq�ɂ߁�\����t�����V�d�N�1c���jV�c� ��}DE�(}ۊ�/��ծ|���oٟ"��GĊ���V�q�I��Fz�=O���#
d&�Uu���,������T�V6�ž��J4��Y��U��3�;\Z�ً.|\��qܚv���1���&�KUm�XC]��"��,��o�\n�9�i����d��_0�| ��p��⚝���,��Հ�
�͌I/��i�d����н�=�%�y��$����o��|Տ�����	����m����J%w!�ْ"�U��=�\6�1&	�����\&�:�����m�s�\73�}~���<����<�B���N���c.����%Q_!��;w���Fjg�S�Ȱ��X, lw��A9�c.O`4@�=���j���j�z�"T[�ޔ���W��$"�ˮ���`�����XG�ܡ�g��^d�7�WmM!i�F�P v2�{��8�>���-�g�Ex�-�(s�b�����"[��	J��9{0��Wk!o��V�Iܔ���Rl��" �G[���D�/����2�!��n���,��Զ;�ٻ���[]xeMq�vHPaR�*�{|���$wq�mw���"ռ�1R6;h)��fc]~���h#	w++J pg�d��2�B�,���\�m�U.,T�F0@��X��Я|���M�S�z�-P�zڲ�2<�����諆����[��ĻܶO�[�m�V�����1�D�~�@'3y���pv}�[J��  l�a�܉�@�0�AX��o���}XGG��xUq�>�u.!��~���7Ǳ�)n�4W1ҧ���/��T��fl���s�|��������i��?#f]YS<�-�fLW�ﳡE��<~p�i�ǋ��[���v�EU��n���Ѧ�W��gi["�1%g$e��txj;�.]�$�B��F�@2Fj�p5�s�/��N�O�U(<CJ#���i~��zl�E���bm��AO"��)y�E��+j��$��c�����=���G����ID�Z3fb�s 3N�0	�MB�N=I��܊!�ּ���>���Ȧ.�N�%ֺt�w9�W�v&U�GGJ
x�[khˉJ|k�Y�7ŵ���[3�����<o��#݆9�O-IņA��R�M.D�9�؄LY9��2A��O���=�2�۔k�ޫ�]y��_�lm]`;7- ���s����%���`��ij)hqn���g�HEy�y�ϫ~~��h��r�dH���t):��������G�1J�:��s��v���\�%�}��/s{���Y��z�]�6�#�{�A�}ݦ��ӫǫ&�r%����C��_����;�.�@DZ��pOSs���5��~Hs�p�]9M�kǍN�6�N�>�N�1��)ꑷ��:0��ౘ[���80�m�-���;�����v�g ǔ;�&Z�cD���f%A��)j#dB�Ě.B��XnLx�\�¸y1B_s����١�>�A�`�i�"�K�1-Ӥ�������v�Q�p�<��6��h�_�b��xYE�c2Kx�\���6Y(2K�-�f��Yؗ����B�J�YR�ٹ��!^[{wԟq��xvt��f�[pC�o��\�6R] �Gf��D�ٞ�,��M�u�Y7�;c�����ic��/C�B���̚V�T�ٔ���/4��Z��؝�F�*��Z������]���K���.��"���wvW�-އ��"L}�8VՆFJ��m%;,:	PE��u:�~�C" )�,,�L�� ���-�����ˇ�Z��\��w`�G�U�����C�Wq߿K���ѧ<�^>���_&Ҹ���ÀS�r��ޛ�d�{�Xf�?����^�+U7������H�u��ɛMONv"�K�xp~��\'�Z;b4OKQF~��ef������F��e�<GE� ���>.�ʢY �t�rG����GPS�9��L���n�G�a�B�k�,�z�ߤ����� �t.�\���m�R�$"Q���%c#p����<ayϨ���v�V�s�cH�I����`Hϡ ,�����.i�J����
SX�ς�����*��K6��H���1T�5dh��x�J{�}��iz��-KjE�4j���P��]�E�ƌ��F��-�0L�00�S�k=����1,�tQ`v`������ș��$|��+����S��/^{����V9궭���_�:o�HWSV�h��>^����|�Q�H���z�9Y�^E���cU�JV�\mQ�ׯ��e��E:+�����Ti�i
_q�Z�1)T�8�`U�ãbBU`q��H�����!A�*��j�o��rR���c���W��_�cb�Em;�d�}V*�K�᯹~��m�v,?T��W.gI�ښoc�\�_��s5�d7 �_�V�rr�[�u�^��R�&�RXjqְ�dA��;m^�*�l��=�T��?C�=��m�0��f1�t5]O�������<M��)��}�^����}��H̧M�������=.�bܹy���o4�+5������-���ˎ�x�O�GH1;/�"������^�Hh�C�AzE"�kv��Ԩs��"���j v�
]Өv�C8�YCf�h��%��J�b{nx������iu'� ��b�Oe�;���}��nD��\��Nll�ul<*3I68ӊ9�]"�j���ĢQ�՞�|2��aAu�2OIM�i�� ���Ж�.1�e��,M�N��/�}�666��^�+����@X�{����Ǐ�FM��n�,��&$@�_݃]�8>�6v�8wn�K�z5aȆ���McK�>�@�3�b2qoHɹ���E�T�f[�Ϧ��:�OqU�i<P��t~�1���łQD�~�lx�鼍,�ٙ��1���fJD`���
F����x��%�RO����Q��*;BB�B�������!���W��xK�4�O����P[:�,XLe�)�_�3�?��������]�j̠l���'�Q���F�5<	ޢ,T>o	u����f5ҊƦ��RE�˫�����u�\k̺�eoq|�wzG�U��{�N��≡����vM�y���޻k�&;]o�(�L�Q�Ӈu�H���u3�������:��������)K)�l~���~�2�X4��B1�#����]�:�gҷ�h���(����}��#��,�8��]�th�g>w��sT��]e�|UvҤ��1�����|*tg��x8�o�T���8�x,�a���Y����E�޶�<Q��9�9\T����MZ�-����QW4	���pCO���w� �1X[����*s��FL�(���H��	K�nV�q�i��]�<|��q&� �\��~���Aʑ}�*<������m,0ן'D]��ʘ�wx�@�P�:W�oW�ŝ�~��!wɉU!Nм��.�P�٨�j Bv��N����|��m�����)�qN�����jZu�������� X�kq�)�Tψ���Cr�A���0�m7=�l�úMf����q���~�vR����¼�M�³�b����g2���t4�hXq�'���Λ��31�"��o�R;�?�ZY���"�9���6|m���ȫXB}�I)|��Wf}t�$�L��g����ǚF4�����c7����4�S�0 j9��dj���teQL,`�=S��P �O�}����2!]��ɉ{��/���n vOޚ�H+����M�'\d������	�߿���v�<�sY��&����c�br���h��]�p�Dq%�vH;��+�P�54��)����q��ŒM��?�/��I-ĉV�SwR[�Q��nSB�4��(]oL�[���ث���e���#�̳]e�t@c�d��UzH�E�Xt0��_�a]4Y���v2��b��e���(ϐ�=�Ǽu�;K�ɽj��й�;��?�9!IW���EH[�*����|���ҩJ��9}��]Sx�*��~�,D��c�R�U�U������X(O�봇&M��ү4�hR^=
5��}}�m:�|4:�����O����n��R(ö��>ԇ0�� �	�GMy���.׽g
Ѓ��w��[��:eo����2�_O�W�>XJ�}��܂t=;���X1�x��D&��E/bѤ(�iZܨ���>k�eo��~��{|7�|JQ��`
�PH鸬n՗��ygo�:d>����c:	>���Ih4�����<���,�根��h_5f�rO��QO�
L�k8i2y)���4E
E��2��?�*�&v,��29�5ęn��ã_�:��YB/���mX��=Y���
���ǹ�T0�%-�C������n��S����Hr8I�%��xgjm��?����f�pCﴆ���&�+[��nIt9LG�惋K�Ejˊ���F"
���r#�+lQ�ZA��'�Dg(�X;wᱪ^޿6�_ԫ���Z����m�_�X�T�2+vp��]�$�$�ه�| ��m�=Z�AUTJT'�A�)4	~U	qA2gk5xD���l%�/�������cu��:�βZ��:5&��V�C#f�H�g���Q��ܷ?�Y��*�����*�����k��t���؆8�'�D�|���[І�y��f6S�� ��cc2#�5�oH9ds�oVI���NZ���ri��5�z{�_�z�ʰ��Iq�h{wC����,�����:d9�p�C�*�2��%���Y��l�������xF�i'i��7 [�4P
�Kc�d���D��w�Kn&_�;y��WBۻP�e��ٙ�:��}=Ou*[�(�=I����Σ���M�Z�B�6g��I�I	M����|�J[�4xs5Uq!���8<��E�zp�;��c ���B�z�ֿ�fAt�#����,W��0UCV?����>OE��9/��������F��?Y�}���o���/drXK��۶�6��a�݇d{��cg�%K���2~�a�c���|�k)���]sI�%~��x�L3�a��*n�\'|
0�
�o8~�WweȜ�nQR�G,S/��Ȟ������xd ��R�ɭHz���C�O����ϐ�WMSlN�j��p����|�c��E���Э6B��h��vs��R	RׅSݐĬ�<=f���.@M݁%��Gp��	���tv~�rݼ)	|$W�Ye�&�f��J�|CR��s8��Q�R唑
k�t��|���Is�zh:��,�
����f�k�?��C�g)v��F��޵5��O-��ռ�����b�X �2�/����Ń�!��/�;�`;�BG�`��JA�����-Gʫ̃E@�����Ao�����[�u�M��vdd�P2e�d6�a����,�{	�ǚ���5;�w��^5��62��ؒj�J�na�1��n{�%�������G�:�=�{���4m$2v�K6.f�J��
�i��K"���k���fs2ym����̩s�^�k�!���t�Fܘ�^��!p'�ᙌ��<p6���H]�f��>��b�˶����d���)�?w�<�Wr����4�Z�E�s�)�4O��Y$C��yg��|e��.�\��������<T�����!��^�MNa 	+���9���`��"�]�(a���5���uV]g�w�{�^�	׏=X>SCs�L��Dk��og<����;�7ѻ�}F4~����TS�&+Dpl�̨-*�����g��������n2�$�JGv��uO��\e�Qȹd�(�I�h���Y�v�	z�qo튿�[|�&���agD������2�5{���R��$ŗ�T�^�v~��E�>��H�}���V�z��z��0�\�"��ojdS�I��|�C3��!����6��)���wu��KӾ�y�~�Q�����������2��.f0�8�Q�%h󖖓�"��0�K�c��$1]��XL��i�8�+l�������n$�]���	θ^���Sw@��̂g��h4+�E��.zW�VQ��gh��o]K����%4iv�紖O�p�|��F��R�֨J3������ǝ"�j1�6�r�Oa~\���s.K-Q!j��������rZ�%�=G(m�#f���.��W*�՛�����V,�_�ʊ�#^"5��:h3�*��Ѣ�$t�<����9)�O��>�G�L�'���Z�얯e� �^��ǚPi�i�~���&J�����<F��UNT)�P9͠[��2�n����#Z�UYΟ5�X��\��[eE������BÀ��~�x�2=4�*�J�-ݚ���Ϊ5��L�%��'Fq���K�{I��cb<q���-n39�+?���놦�R��X���=�;z�ɫue�n��]?��(�I�cMmƾ�K�]�d]�����!4b�rs ��h���sP�X��֛* �K�Hrs�?�\�TjCe�d �����\ϭ�j6�J*,�KC*2�p�GOj�Ўxww��y5
�
�������v�	:�T[䎆���p�U��\DJ�/�*ҸoY�������c3�r4�t+���#B}���l��R�:��%Zʵ؞?M�
�����~����f ^�!Z?Ud�q�Ћ�>��z�Q�����e�+��{���KGt������C�w6�?�b�^}�l}>9��8����!;����+��<��e�,-*A<+//g�}����J���Jhۭ_��(�~�O�*�!%��l����`9���^��\�<KV�5���#�;�z���{��ѯ�O��9]2]4_��0D(�T���ܻk,uqQ�W:�v�PP6}�F�$ga�TS���3���a�7pQe��lW!�W�v��F�R&��|�u]
X��4w�]�M��?,�1VW�;�	{��?�E�J%��C��h����k���?��_���Ű�~�R��	�XN��4�z?;����������Rz"d�ep,�7���I�;3zg�.@�8Ut���gl��=�C,T��%���>�V��l0�D:� �H&�+� n������A����٨<��hHd,L���`�A�(�C=}��$=Ţ
��@=�@�'�y  ��E�u���;��)ǚɧ��i]�R1��]��㘚=%w�u�O{{W�b}�:��Ѧ~vw�!��N�&�[b@?����$���	؉�8�X}�"$�S�`O���8m�w�	������vyaȮ���+�P�����ڦ0�4:�n����ߘ8����>�FXEΔ�4���{Pt\�*2}aq#�3A\`�/�!}�o=�ԇ�Ec�f�LWw�OW�<
����3֑��M]̔M��[�X��OZWq9�ٹ((-���VKU�Ɓ��Z���y�M�:������P��z�����W����wO(�[��׻Y��BC����pٙ���|9]W8��^�Ȝ�n~^�C��4����C+_���NLm8��#'��f�^�6�|�܃SB�g9�}5���x�s1�)���u+�et�|��e�9��·�WP[ѷ�Bξ�l�.D
q�o�Q��bٱ��qΖ�E8�#�/�gJ�!선�s��%�;��॒��7ۻ�wg��y~/���mO�}��ɣ�� e5�j�vY�5���P�*��3A>1�خQ��|������B����Y���8q�ȚHa�Zm�w�o��:��Wt���/rsf�#]Y��h�H�����Kɘ٬�mWT�gZ�����]9���M.pd�m�1"�M G0�\�TkMI��7�1ū�������2�����92�^���l��m���G�~3�sYU*X�*�����s�I	#�s F��S���V�9<&�����okZN�>ǟ2��������eꗫ�;J|	�o�H�ϑ�<va�0���W$��ٺ��G@_ ��7mI@�_�U;�����r�[����?T؜a򢔯i0=:��/a���o�G��=�ʹ�)A��_�58G��X�׆�
n,9af�ч�Im-�*��չ+U߫(����vįnGC�T&��0"��Tc������ȷm��O��Dw���5�`e��v�h�������:�Q��5>-
���73ݤ9�/�Ϣ�?�Ѡ�U��N�w$����N����֥Eݛ���I��:�<��~�oX�nn2�'���b���TCQ�:DM�\����]%�d�iw�����9=N(OSi���kʅyY325C���Y�j��d8]<� ���P(��$,��B<s{�t��t�Qj����u'�S��W&�5S��[-��5W���A�������{��񛴯�����ϥ�!�>��=��W���}��}A�B������i,�#�aJNk����ܞ�:�HR�O�
~�L�.��n��ח8@�H<�� f�����W��Pѷ����:��Q1�õ��xi�{��<��8�8�u<�ť�.�x��W�m1�Ӕs6D0^�s�O�-����ZMf�ą�w63��:J�g�v�2��'\�z��z{�XԸ�I��z�IJ~��Z�q�nd�]��VJ3���Ȏ"�n�;s΄�<S�i.��]>kG�'��F���&��뵸J?0����θ��QM�!��=�9�����ɛ�A9������p~q놸ص��Ą��YzPX�9������X�m,՞���A0ֺ��kU�'�ZV��!�-WΓ����������:����]�¹�3��T���T�ѳ2�'*!��E�=#�%1	q������Eim�gL2�Tn��-�t�d�Q�E8��b�$+�B�����+�j'�o4^��y�%P���u�����z^˽����)��n�^���fԄ|�q��_�l�w|\��^��_�)&��ȍ��%(�ZȄ��5Q`��8	��7�>�k���J�����n��ޝ�ҿy��N<@��±���lC�� �V<>/#:���R�S(�R)����D`�^�O|��5;��w�c`��!(
@��
���do�)i�+��ܭ>S46�!	�uP�l�u
�>��:ާ���st��I{*y��@[�^����g���칡V�gR!��3�yUņ!��7M���H�>0ԏ��an`�h@�	ѻ��O���Y�8p"�.�z�5	�ԝ�ʱ
��Ƭ5��SJ�d�?���)i�@��R���F}'�����K.ń�#T�G�\��:Хb��$r֓���z�I������#���/KrdҞ�ԺWI�A3?����LPV(lڂ�����:��l��%O~�cF2t>�į<��O-\{μ��^Ƚ����zL�j���N��:?⌣���0:�%-_%�zdX��=�wM�ۻ6e5���zr���I�l~Q������Oji�D+ڲ���ȇ�����@�`X���"k���qi�5���+č����]b���T�EK�ɬ�H��k�j޽�,�ݡ�Wڏ��Km�J�������o �^ɜO��^�3����C1��V�
��?T��&5_}�m�}�����J��͑;C@�?�{��`o�J�/+�+q\�b�� �\�:6L��f}����bk�Gg��p�G ,�ދxa�L]�
`!��{.���\�O�]<����l��u�O.�l �0�&@n�'�zu@U��1���kw��v�a��{\���MZJ"js)�4 ���o�.v�V|�]u���7�1�7�����g_��#�֌՘�U�9�z�\z��zV�~��K��_�<50������b��%�4�M�^���������O�Ϳfz÷��^��!����rBm��FX�j�"Hxt�%����\�g������W]T3	S�k)�C��ׂ)1�V���[�m�x0X0Ho��.[v�4l�=,lg-1�@�ykqd<��ʟ�¢3a�:{z�b�쿡7���'Ƹ
W7����{5l�y5&s�0�;z@vŪ��$����y�kV�Z�O�t6`3���%.��G�<X�J�^��f}��J��g��mW1I2A��y���BȆ�OS�.��t�{�ȍ�ʫ�|��A�����Yi��ԑ/{�`�
Hۄ7����Z��2���B�n>�Ih���o���mR�k�������?/7�'S�5П�F��5J}k�u=�ɾ���9�����-���i�$�/�l�1�w|����(p&w���7���㴲�bY�+��t5�r@�\f���N?gqMs�B��P��ض[�w#a�Q���R�ǂ>[fWR��~"�d�8[�9@O�g�S��'��#O_\�1���HW	�^�/ҙ��5C~�ܺ���;����\��"}��l���@���}��/��)���sy����������k�����!�ǔ�)�hK���ҡ
��0�V4���dР�؆$D�
A9 ��p��HҠ)���:l0�]���uέr����c�q�N�j�0�0�}qA��ϱ���.�4�A�n���� �>�+X�R(w���5P�.��'���5E+�u��w�z���;l/B�mM�V��a�[�g���H�Τ呂%���s4���{�c��i�f��������uŢ�df$�ѫg8�6����g��{7�
��|�OBV�c���'1#�A,ց���D��c��ʬ���椅DNke��籨t����I��]8g��j}�����Pwp=��,�����-��O�����9;y��h�2�7���<C�>p�P��>$PAH�-b�'/찋���:�2��a�z�׎��pA�cd*��\�Vy�P�b7�[������@�F��J.*X�r�.0���~/�1�u}TРi1��G�q��C����:;��3��.{l��<q���ϼ��K	P4���.z�:l�~�g�����3�d)�+⭓`�ȉh����DO�sh
�l�풛?�
Elw�(%�{g�;�e��z�6��o6~�!>o��DW� �8��+�29(����D�{��zF����>wawJ��e��j�����?�fj��"n�g� �GJ��m�!�$���|�n�]t��mO�X2,���w[ᡔm�h��䲩K,�8B?ntϼx)��7uX?r��a����$��=v:l�5 n��;<�n�N������_Z��^��`l�����]�X�;�8��E^��Z*�$cu�r=db�C��ݮ�[i1����8���dn�N$_ �u���Q�4ڒ���@�-/�w��y��%[Q
�*eL��u�
Yxa���b�tM�ZC��ru���w���d��A�ϫ�ͦ���]��;�!V3�bF��ȫ}]��d�C+����O�wo""��,�-$*A����\_��^��l�L]	R?k�	@,�.�cl<��Ҷ�i�-��bD���k��ͫ�TM�����g����2V.~1������FڇvzfN�v����
��U�-��O^8/�p�ڰ����sz*x����FW'��2@���m?�����=���խ�z�)�DRN�(s�+�2��*_F�
	Ag\�f�LU���9K_�e'켣a�:b��zs�y�ĭ9�E���Q�Ö����	�-���&���
��S`�N ��jb+]W�e��m}f��kj�K��صl����vo�ji�[�rx5
R5���}��fKԇ�����ȯ3�y��c����b/S	��C�"݇!,_�4f����WK���Z�/�:(��dg���U#QB�3�{���oL�7�L̡�8��KCH �@�)	��(��s�kPh��)�d"��-py�8�&j�8��8
��b	�do`�6,{1�K�.�T?Z)@UDO�\6�T�+6#4@a�衢����N��E��UҊcl�nk�&_�n7���z=� �dM�����ʎ_�ѐ�bRw��������C��4��-[1���f���\�5�a�[�U� �=� �#2����םU��Z���.���#^�L��EF���X~�~��e>�X5��['�<���iz�C?hK냋=د�c% !�U�b�#s~~)�6�/�v�y�f�;�$��Q��~+�G�
~v�.}|hEEMx�Hk�EG�#3��=g�3�g��c��'��B��xT���˦��ќ;����hVI2��N�K�����̟{*7���[LY��;���P
i_��U4�F��H��e�l\� ��@!N���mr��v�2<(��5�R��b�Z�o_�1��iy��b
*�4"�:!V��]��9����Cl>y��Z��y�vF��Xkȡ�شFp��OL�vi���x��m�\|�qwt�P|�Z����ܮ�`��Q��G~J�M��5�D(,ER;���_��DY�}蚐��CJF���B�x��}��5���%Sf�}	 ������n��G�=�)�F=
6��)�nW�ǥڐ��%�,R�"/{��}�j4b�W!�J�"���E�b�	��ū]w��3�@��2�B�SA�c�e��?�
r��R���;������)�e�x����l&j�:��f��OTY\gߙJ�DM�/�U�Zz��C�)�v����J�+�]	1�i����>�r 䮯W�7�m{I�iV�fۑt��ל:�������Y�%�Ǚ`������ꍍ	����CPxln%L�F=%7��Ql�iv˵u�B�@EfK��rg�x7*�w������wHx�2�d�t�xW��v�=�y�zY�g,��'�M#Rzyf]��pJ�qt��Cs����w0��}ȁNŴe�y��O֡��R쓠�g����TF���j����͢{��[�o�٥�|Wf�K߭�O�#����;���;�-{�7&�Axn�]ҫ�ą�J0N�4zH-�J�>�n,�W�>r-c���(�hs��ɒ�G���Ɯ�H٥�ԑ�=�2�g�mT2uF���,�9T��5פ�q}ī�B�R��UTR�8ap�3R�@
g ����m�\�65�����6e�E~��s��:V5mҤK�A���E�X��/}���cd��l�ds�d����R[�N}:q1���nPށ�2�D1�����=lai5��}��萨�vdTzb�Zp�¥�B��e���}���xA=��:�J�����M�د�#9��������}:P:�8^����C��������-�
X�jf^J5��/��BE�/X3DԪQw`{����_,Sdp�K�_�1ϳ��?p�܈�x��p.6E�̬~T�y��4bǯ��$���K�+����:�{����
Y���<vj֣n��Fp��U��!',"[��5,���RѼh�C�΅ی�{k�l'̆R�GZ0�h��<M ܎���G$H����a֮ɪVEg��)��_Ι��|��ۻ2l��y4)־GU;/_k�h�ߣ�@a�H{��p��0�&�e��%��H��O�kL���
��hx�G�0��dB(*[�SW�Os��]��U���Li�d��T��&��(H�)�x���>qzT��m�2�X�)1{����rбP�߶��3߬~7��~@9=R�'׼�/�6��r2`�%�vϸحԊ3lX�CA*�(`V���þ�(���~�ބ�������	�:��]#��eo����#�.ŀl����y���jɬ{� �CA	棻]�B�K��E!Q��O=�Sȓ�^�rYD v�r'g�K�o �6۴3Q�4~����u-���&3���\k�b̢(���L\�d\MT���?ף�x���҅
G�3�D����?
�?2��w��Q�f����Z�3<M�7�ǑW^e��ӤȥiJ�O�_�\��>/��P�����B�4=z�m�V��lH�RJ�	$�\����b��t@�z��+	>��m�l�>�1��q�Q 6�ZY�L��<<O��c�T��+�k�u��֊0�J�t>\�����������j�cMk��!)��a'�����p��^���W��>ZH�^W�a�\N�����鸈�	C.;u���?~�e�.�:��b��(uY=���y#u���UX�]�ÇK�vt|�0�eᡆ��?3�"MA<2n؆M)Ȧ��%U�Ԣ&�	�S�Z�����w�dͿp���5�a�_Y�Y���j<���#��	�zH*�*�	�x�(3���4>�usmr�ce��,}6^��E�����9�OG��������T�V~�����e��8s��p��;���@�̎�p��>��j��{ts=~hs���J?&|����L}u�R"(T"x���G
�����2Nʷ��H5�rv�R�g�WK�}�u���η��A�{�C����}��0����F�u�Z�g� Ԯ\��Hj^�A�.U+듮nϿ��������n<㣯�K��4�W_����b��؇�����'	�V����x��E���!X�]۰��D���W��h�<Z��t!3:��|���jES,�Zx'�v71Ի?����r��zg����OGZU~�����y1��7>B&ĲO��2��d���-�����>�B�Ǜ�'*|Z��,&������_R���(�����9�n)�������+���nOc��Y��f�d$�ɀ:6(����p���z�]����Z�0gnuH�J@`�����#٣x����^����b��yS�ݴq��^S+��5�Y}�U�Y����w���o�㼹��U4���un?';(Qz���}8c���
@�ڳ�����Մe������G����A{	gjӁ�'�����G�y���Yx���1p�"����̴���K�i���*}�iZ�g�U���?�����*B�/U�>��CK�x@j��l��*1:�a9i�ǉ{��J� ���m�����D]OG�~�922�6�Bjm�O� �X�SYl��0���dp�
PΜ�)���{i��	g�FZ��7�89�]�Q��=_�������P\nA?TJ�ٹ�j]�'<�.R��70���O5U/PnzۍTV���٥7\}_��yы����L~ش���T�t�r��Թ���3�C*ȯC�ƛ�gN��!�����)��9�2`�ia���{	�:�B_7�?8�;�w�3��~�8�my�����z�����'S����S���Xy��k�8��R�9+��f�R�!��[a�xZ�����e�&vy�J'mx�}wP�������LTb�a9��c|����|N��$�ߍ�<f7��@�yrL�o���쾨��ݛ�9!����^o�r�u��Whis���D���}���t�_�p;1��u����J�S�z���mˎ��N�T���&qt��Ƀ�	7:˕9��������X�F	f�6�R{�ۻ<�ּ�#��3da���d�Wst~�s0s�v,7@<�����z������l�T��\!B�9�7���o����V�\q MQ�5u
l�^g�<���v���!�S�֠���?��eN1�e���.l��@i�<���!�s��Xl��������ئ�������{Y��5��)P�h"��~r��6}�|�1g\��YL����IߩG�EM�3��E�v����&�]���#>��z �f$d������~����Y��i���|���n��܌VIS�62_����'+�~��j��Ozꙣ��Ӭu�¤{�u@����aX����R��ib�mwHF�2Qu
�q�o�R�,\ЋW⁭m���u�8����]i<(�]�q�VĩD��YNS��, ���(x��)��8�{�W9��s�j�,��#��cŋI:%�}��⚄�8�VO"!RaVRH�x3��/��J-��*mj���'?���thAC�ՙ���K�e�섕�|?z⁐J�/M��L���e�^�-F0�<w%��W�$�d���Iz1�Uٗآ�ʹ���^Q[���#�@k.e@c���pt�x
f��~�-���H$�ժ�g=d���)�R�S,�n�Ln=���n��4N/(����Ϭ'�}o&��n�+!4��	1����B2>� %�5��&3@�fBVV�����p�.m�<�g���2�	��RQ�!��RJ�"�V0�M���E�԰�D+I�#I��Nf��NWtIZF���kr�2��z}B�N5���̈́#5. Q����a<e�����l<3@�D����p[d(ma����xÑR�ߖ~x���^c�z	,:�������YG�Z��������2�9�Egy�ݾ�J�q�����<�5��/V�bU)���E�s��Mj*ns��6;{��y�J�.׫�k.����1X��bt�N7)@�����5�F�d4���8eb������j��{]�0����gY���[�xsW�}:��4�MЈVYo���ϥc��P������.ұ]t�^8�V4pꔺ=k��>߅����eT��H��;#ΗW��?�����?dsvO}���QF>������"���^�����*�1�����le��a�̵,�3�	�kY��k�b1�6��VU�H(pߞ����ּ���w�F�U�Jg^����ъ����qso�9� ����p�ă����s;K5g#�S�3�}���� �X�$58��ҴW������鷒�  @߿@�߭@����W#sWߙ�v��O��6<�!���w�yk�N�v�~|���1y���4�?<~8�u\۹��Ф��f�g�5��pu	?�╿ɛ���k�U<f�J�,�\[�����]Fp�?z*6���[^���o����K^�]^����=pK�V���f�i�N�h�t>͡>��Ë�z�NF���\�R?�t�,��|1����,���;|�4l�U�J�� �1�XF�����?K���j��G�(�� �7)r{�y��oKgq�_��(��ҽ?$�sla+|�edV�	g�?���.^a����x�np�f��8K����S���ֽ���N�����t.S^����!�W�o���4O���i|6'��t�Q���F��q����x��:�tOK�tX8���\��#�:e�����d�R.���ԧt��L�d�������]n������7z�6��*V�ԗ������
��ܛ��\�������޵!��{�)�څ����ׯ0�^�W�^��> �%���f~����?��?O�7�����f�������Vl�*9/�%��`.3����\�16�!5��E�Ѵ���O��E:S��>�jF7�o�r�>u��$�m�F>�J����8z&���(��.Oa*O����A%'ft|\�?���Vd߅B�M�x����2X�(��XL�Q�F��>?|��ׇ���������?:���ɇ]�'��L��� �kz�y�.�<���[r�|�g�͸��~�ǖ�p�h�&l��A��v�]L8T>&~�=⭸i�R��J��Y�ާ	Sx[�t4�d�u=aK���?�����?�χ?���U*J�|��O��O����놄҇�2����)��3W�N�]9-����	y��Ü���Z�Z���Z���fw�N��wE��[!�oܫ�&m!i���.^��^�#?��<ȝ���F�K9�D�g�@�J>vUH9}��u���E� I˽t����#44*:�m���)4�拠n$���Ъ��z3��4�zx+����g x/g��G�u��W��Ꮧ۷�L'[��5�eVNt�y�U�|w`����_����y7tq�x䒎�J^G}��tP�PYG�̟x_|��(�'C�^|�����.��5! FG�t[g���M3R��<�~��Efq�C�uD�i�}������`�Eo�!�#��&����O\a��Gnߵ�~8��]0�������;��Ç[���޽3���7�����o�;\:>t/�@~ݻ����ё��=x��o�?:S�z�����(O4M���6��Eg�U>����G=Վ�+�V��SV����s�����W���~2d�9�'9$~��t�  ��+����^���y�.����7َ룧p�A��.ΓlYq�U\�0C'����9Y�ŏ��[~���..�=x�W8�y�AS>io�q���5���'�.��8�_���?w�Y��%<�k�W����yz���t(��<x�~n0C7��������G������d�����C�Տt��;Z�,����-i�+�τۤyl��6�+�ѩ��і��/l]�B>lg0�4Gc��<�Vڭ��n�J������;}E�cC�7�%�	���C�	Ź۠����xl�����p���
VB�Ce�9іG�dr���s����#��	��-3e�J��u�A~�3��/%px7�@ö3���A���o�?���/8��f�����M��t��`��g6xt�Ş:�n%���dD4�^L�8�z�y���2Ǹ��nI\�>|-�йD$*NSr(����?��Up��ŗQR�Z��V�3B	��܆<��xXdd�d�����R�
�R��w�"����b����ߓm���É8H1Lg/��Do>M�{�3?y�����~������u;3������g ����~���|z��ٶc��:/p��e*�W���H����:���D�g���+����m
c�Zg��+��3Oz�̿��1�uy�=�l:�뼆p0ᓧk�|�p�n��;ekaf{�k��I��_��_�L��(t:+$���	�*��7��.?s;@��晫i�_������?����o����~~S�\�ͪ���~������O"�k�����)lf�ra�����!0��@�Dt����v��������P������E�<������9�_B3 e�?3	���oU�K��T�
:ySa�-�5�X���qQ��^pa��F�Ow�g���>�z=��S?2�wҩwY&I#���LA�}#�R�xh�tZ^䃍f��fy��*��s2���.gP�4_�������ຝ���ᳯϟ|ux'���r�t*iT�ߺ�V�Ϳ �iXTVw�θ��o�Y�b,�?�	�)\���w.��|	�����@�wariv�H�=�;8 W!�	Wߺ�1�}|�p��w�,��!=��N.ޙ�5eF#q;:v3r�:2���tЯ��H;twB_>L�t=v%���W�{���nf�s9��WI��B*V�hP_ތ��<�o�<n�yd��ݷ�:���{����*�ċ��O#?�B0���K�3�:�מYIY3�:�Xy�:�[�$�q-�{-��rx9��\ʍsM�3���Qd}qx�-��L�����ԕ���Y�.2�#��e��1�� �~޻���
{��{�G_��ˣ���0��O>�����ٳ�9��<}����3�λ��Ǚ�ҙ����H��Ɂ�F�7�f�m�7��4�]�*���ʠ9e ��[L����7�1 x��ї9�%���]?���{{w�EG�N����ᗿ�U�(|�ⳭP==3��rp�w���lEIyd��M�9>�Q_E�)��StR����W�������;�7�=�w�#�~�[�C8>����-(�?����ݐw�ꬰ������Xco�������4�5�c&��z������	�mf�m{p�$��)O�V���v�ҡ]e���O���7O���L���W��t�W&�e`��*Y��5�u++>��4�w��0�3�%l*�Ȇ��(�<M���D�,��VS3��/^dr'���ї%��͟�)w|��EV���r��;ã��kZg�q��F������_>��g����V�3�l�҇�=˭)����>¿o,I����:�겛�����ӟ��ѕ_���W9��f{���]e{�x�^K~��w�ڹi�F~����O�?������㫂�3Rp�O]���t��w����xڜ��\��.[�;���9��4"����Ow�E���S�_e��M�e)OsN��[���ƒ�\�U�i+8Y\ھ�-=�*l/+g]��}�=���S����Z�����?�<}�+���/��?~�ɗ��׳*�>BT,��3Y���?��?x��×�����_��t��>���мȍ�_%n��v�so��W��Y�����\F������s+h�{/�_)��[��17%F�}�-��,�?��JHL�>�M 	z��{S1�
�+� J�  �f� �O7��O����i�[#*����,Yv��~�0��G��=O����;�o�����έ�_���=��/����_���I�|�Y��}��\%���4�7��$�u�*��r�BAy���m3���x~��s:�f߰&3Ep߉�W4h�I{Jb�R���f����T�,.��5����ʒH'#���g��{٧�x�^yM�r�/�:���Ng�L�����_t�$Oǣ�1iH>	{yhdV��U,.nch�޼����w�x؛�����O��S�{����Oi��k��y�qP�f ��P��V_Y�13㪲��d�`Tcu�A����@�˖i!3���e�����i4�fM>�藯�?������탍o��@=��P�J��̢��ʌ���w�~/�v��R�ߙ�k齙
��H��˃4b�� "�̍9����)Ne�2��Ƀ��ߍfk �b�u����Y��t�_u�3:���m�����t��d.[Hg\�ܞ�����I�4�&B�ҭ�[��e�Aٴ�`�� ����0��uː��/�� ��#���Id�������;z��dK��g_}u-+#_�Ap�WRv�����%�� e���3�{���Rѕ�"�]��u���t��~��&���	���wr�>�(G�ep�#���7ۄ~���F>��Fh 3Öt�N=h6Ί���t�@���n{�����G����e������F�x�G��7k���t�����jWԩ2���V��d�,���}�����o=Zh���?n8f/����;��N�Ėa�#��c����r-̻��.<�S��:�_F��ˀ >���q��=��?�4��Ig�7Z�V�Y��s/���U�y�S��`���qG��<l��#�>����_{���|Kܚ�S;���Qވ_��ɯa���8}/~��-���`�������`���K{�YyQx�|&ũ�OYfÁ7f��4���-z���?�B%�*~���Ħ.�����eWL*������̮O=>�RGө>��_��<�և�����J���ve@'��5�^��6�x���9��,+6�Hfd_��ܵtb?�çIGv�|�մ1⡱��2�A|����<C���V$ա���������{/S7����_���I���mb=g����9<��v� �m����$|=�������E�r�l�4���<~�`�������v����^��Ι�o�����Ç��y;�_�֮�������9+�v/i	ogE�\?|��=�����=;���{���O2@��窃��7��͑����o�����b����ﳝ��������O~���3lP]��t�(��̡���*�q%�de�����lq��Ș*[�t�� �x��R`L$���������0�
�p+,k��n��E2ӫ�� 
����&���;��~���}�Gӡ���P���I����f�zfG(tȞ=Y�5~F�����������ï��I��+�~q���t�\��� �oo����CY�ǰ
(G���tw��ZaDyȹ��@^+�I��)��,�.O�U���ǔ� 7��قx�o�QVZ6#�����"��u�LGL�2���گ�4�Y��mk��I�F~)H���Hsh��Ӳ��<�{aVYn�����n��C�.ȅ���������ܹ�ӱ'�T�V�l͘"��2��f1�@S��4#��5j�m�('e�5���t��G7��t,��L,���Zay��8�cU�I*W���۷̖g	>���ҁ|z�d����)O�-ن����܎3m7���g�,�����3�k��&f����:������9[�n�"��̐�bN��
�Nod�{�	<N�
?VqF��K�?��3(�*�w�o���b�G��Q*�K�ӱO��,]~���F�\�t� }�+�52&&tޞ����ε�f�5��Ɨ�1uq����ﶩ4�z��&'n�T�W9ǯ
Q����nz�<C��S�O[{�W>�H}��ש���@�������7q��zΕ�͹��{�-�_��Q��鋬�$�#�t��0��f�4��f> �$}S�J���T�ÓU�W�x��Z9Zg=�Í�1�n�q��XJ�ߤ�E.7���O���zy�$+4�w7�$��@���G�y��I�ĝ���y��6זkv��O��L�����U����� �3�E��0p�Z�c_eE��
��hq�{����0I���R�'~��.l�����������,ۏI��gBd��8���-��k�c�"�F�~�K�,k��4�w�L�0��)��U���)cڬ�t	IQ?��5EyҰp�0�������p��#�(���'����
����q)���]M��Y&Q��&3�8L���x=`+~q�C��C���Hu.�I�U�����͉��UQ����'=�]Z��OF��W���o�[=dF<}n��e+<>˪{�a������-f&�&5���u헳+F�4fV�7}���n���O[>���3����j�ץ_���<�s ��Ip�����Z:�O�-VZf*�aҪ���H>�Ԗ��<��_~�m���5�9�+Ϸ�T�/.=>|��7����_����n��p��q>�l˴�O�?>�Ar�Z�}���.�w���pq��û�}o������ô	/����P��:l[�|�ˎ���_����Y��,��&��'���b�9y?���]v2���a~eD3] 7�{��w�������$x	Ib�PR��G�
me�A�)ӅGj��O���+����I�H�����C[}�L٦���H1��=�*�48: ��y�T�Q��%�;�lԞ**��9Ě�Zv+n�J��� {�uNe��+�wogV 
|5�w3���%sR}� �w�xꔸPu
J:
��O���;��Lj��>H��ay�۪���Z�B��^~:�`�ڳ�V#������`�Ϣ�Mf5��@���/��Cg����Xu�,�
�4|fT7��o����$��=M��<���g[����^���&��}�32�����W����6N*�/ә��mO:�`�$�D&ԛޘ�U!�����0��7[#��*�'�F4�_��L��Q�%�����۾�mA�s+�����~r�Y*�_��㙑�O�O9�~����{��=�V�~�g�,���Y�X~�T�f�L޹�^:�)_d>�-#Ɠ�7KUq�2ϵ����	���̳ ��D��X�Nq�6�"���G�"WyN�2tth�%��>�����7Z���J��y�&d�f�g@����=I�;yf �C�㮆�m�B�wa�Zg>2!o��"�v�5곧�e��t���������4�h��D/t�-/�S�ԍ:�.`�FGt��ŪO��NDFf�E�w�aǯ��q���ԣ�R��z��If���Y����K�yiF�Af��a�Äʔ/�4��6��߽�n�أW�1�Թ��J�z��/ENh���i��N�t��_e�I�Y�X7��؞�&,��wj3�%�+Xn�j��?��dfE�q�&����/���a�\|���e{��5��~���a��n�,)��F ���NZ���u�q����ȎN�1��W�h2�����3�sؾ�6�ބk�0��]<�vӳ�/����sw����_�՟[<ֽ�_[ع��^���=~��a0���<�+nn�X���5N��fglupa�މ^1����:��3}��v`����B����4�� �KK8��iN0�Ѣ�V&�4|�
rJ���.��I�A��I6��������'U���G\�!�k`�<2?�;6/�`&�_�+�5�Ң���pJXuM[u"�y9�Aʓ�]�duw��W�ڪ����2�x?+��"��������g�V^��`3h�=p����T�3T:�V�ѽ�:=)�E����������~���剟m���ͮG	#����L6�!����oo�L�����i���z�a��o���`]i���3X�3�{ٶ~+i�C�����~��lmM�f�a�B�+iB���'�7g>l�R/"�<'�4�fфWy:�.��k��`o�f�Dg��ZB_�����-y;�����:w�_y�A�BD��b�Fi��2�:�Na҈���dnD0qG�_D���҈��t����ύ4��}7#�{鰽�A��r��͒�=���<�&���3ڝ�FʨD.f#�4��V$��}={�Ʌ�kX*#�Q���8K��U�(�C[Ky*"a*.|(��%�� Y�&��¼*C|�
s�}��U��j6%�A�5�9;��,��Ӗn�a�óh-�~��-�8�?����&!	=2����n?�E����>Laf�W2:�.|���h�l�ӱ��A��f��
��+^�����tʢ�#����\����{��efn������i�@�`^� C�u���2tv��ן�d6�������̻��������Y���������[9���TB��t.�Y}�s3�=��u�}�������̢��e�l�M�5F�/���AF~���97��ieKQD�� ��h��G�Τ
*���סe�|��%[�1�2C�*[�N'�a�6�ӫ
��{�=9Lf���v&���Y���G�fk̐������ՑIV2�{�b�T�z�\#��y�<�"� ��4�Z��?{o�l�q���������;@PԈ3�F�
)
��Y�����7����ٲ(�s�}_4���{����̓���hE������;�Ԛ������U�)�ʊ=�X�a�7��F��O�5�(��s�u��m3`m`W-�(�O����E�ҼP:��\��pif��ʟyj��7��Ҧ�tM4�`���ӡ-�U'+N�l'���)Wy\��s�a��B�>5�
i��,�d� ��U W�m��:PQ�
\�u 5�l9�G�Ե� �/r��1ɩ���L�����h�K���t�OZ�.�G[[�?�80<i��p�_��ƫt�0���myk�Z�tbnߩrm7zڗ��t�e:��z<Yr���,���xUN�]i�ٍ�����~���w=�K7}ի�i����t#��
���5��'0�u��`���م�x~���W7�v+'��ۤE�.h��*��ҡ�|/��򎾄����� WphVe���	�Vr����	�#|3�^�3�5����}e�F��Қ�.\���d�p���\��u��/J8�����G*����ӿp^}���/�Ŀ��T5�_�1ƕП45� ���8v\p��׎xCc;9g{���J���A�E�W�f���`�*7���>���c|�Q�1A�'�?�P�j`r|M�2�%�VU�7O]L��[��of8�nܾ��^�I�G�E�c4 �<T�
,�
��n�ob��I��H@���(h�q��7�<|�/6��0�jb~)V8��n�:Ǝ���l!VI�P��;ws�E��ulx���>a�X~�<�R�X)Lm]rl�~�W�:��!LYQ��)�lc�����.�G�������P�
�o$����������8m��6�["��T$B*��a�?3�n�]�SK�N��N!^g[G1�@23'6�Ado�&5�)�V�/�K6lZ���I�?M�q���w�&���(�g-ũe�4�qdL�hue�����,[����Y?�O�)����tơ@��Z���+M߯^ڧ��Ӛ����P�Ţ*�֋��ՂHX��ħ0�Ū�V�G� ,6���˚cE���햗�ல��껞4*!�oj�%�e�ݼ�C�_��g�w8���շO�ب�j��Ofۋ#��<��+/̉�t.�{з��ܖXQszV{�k�!�y�w���6�l�,��pF���1�f�M3h/:u�9w�x,e������@l�h%���g�E��i�c���ˬ��B'�NR����bz��_aZ��*��+��7�f�8��=;��V��-V7n��&� bc6O)����v��A���8S����vJk��3Qp�� �Dr�
����8�D�ˠ��$-}�<~2a_fY��kި�����8��(�-�}a�I^�y��*��	�&H��uWS��+�L<t�%�r<چ%��Sv��f^�^z�J�=T��d��ٌG�j�|��N�&��p��F��������0��t�)6�mň*�[p'�M�P9ΉW����X����1&zГ�1��E��	�cy���q�%���h� ��$����X�?ɉ̮�Mcȼ�lB/���a
�/qg���Ӷ��}J?�t'i
�W�e��ج�e�?�(g}�<�w��:������;Q 3�
���a�5�����V'�~�a�_S���JQ�@ZV���V��4?�}�w��Sq+�����Jo|]7N��s8���>tE'�1�'��ԩ��P�~�ޟ�i�?�'�OqZ��o��g�W����
/?���Y�~믟��Εd˯p�*g��K���w�+��!�h�c\��+�*'ܰ����$��4{�]�Ą�rs�4B$'�-���R�e(��m-��jB?��Ğh���A�)ɯ�u:�8s�LXS�2�rU��>��i�e��Q>i+�y�^�q �y���I?q�u�����)��9��CHo͛ a(�G���~;���70���d.�֎�=4�pq�1<�>}�ffX��G!L����s����l���w���fy��C�`R�)QN��5�s�C���F�Z^]g��w1.���on�w%߉ȝ[˜Ⱦ��L�2�M�=V��Hw�u:R�w��ٸ�m����uo��N�������Ľ�l�ͣ��s�U���N�)�K�-���FH�jL++���uk�O��t�����d��.%F�e�_�w�B��	=9`�T�����D�.q�A���|��IlpC��>:�\?��(�ٯǳAct&�Bc�\��w��\�܎���s̖c��(cvB؂@Ќ! %у|&H#���b�Q���l�R۠��u�s+�a��g�L���Ky��v�:�y�x�zn|'j���;񺰙.K�-���3�ɟ�:��fډA��3��Z��!@S���4󅿓�XE�b��qZ��_a�	M����pW����͒��jR��t�*��ʯM��3�[�U��q���0��W�T<{�l��	F2�h�:N=]�+x��!���AO���ഉ텭��`0<o@�!D��i:�P�ʘ�,a�9��zlm7U�G#r��Ο=�p�W9Mm�B���f]�R���Gņ�I�f�
>����U:��oN�\�vއ*�z�h�����Cs��=���ɥ�\�0�Bս����:}���s����O�wn��`��xй�
-�}7a�b�"���$��F'Us��I��@���<�]e�����T����_v#c�.�FN;��ؠ�)��sϰʤ���iײ8eJ��AI���T.�g�gX~K� �8�ɥ�mLS��MV3z����,6A��.h�h5\'i_���4�Օ;�{�+L�D6X�&�Cv�h�x��a����[q��(+W:q<�����3a�;�B!}B)F�I�M�(i����07M[FiP���&T��J�0lr�刴8��-Ͼ�^Kaa;�k����z�H�7�)�y/h���IUs.�T�綘�H[�P���:]we-�%>��w㘟���|ͧ\�ex�c��~��#�T\ηZM�9M;��7˲ݍ�wLhHg�/f�UY��r�p��p�f|����W~�a��d1���q���/x#*N�尪�t�Ϸ�d�����S�)�~9��*�g��3a���ᾛvX�4~�Si��շ�îҚ��(Υ�a�K��L�����)l-��D�%/�t!��	K��[V9�/%��V��>ʟ&s��� �iN��pW�]ٜ�OL!/u�<����F]�a���{�m��
G���
<����}G����>����[�b�"خ
��YB�O�/�6�T)�*�("g}��ߟ4�S��s�z�8�#��|^�Jq�"I�vy�3a��<PÓ����¾<�y��rL��9��8�F!7�1�'�N7w�����v����O����(�"O"�O�m-���=��59�<���T��v�qO�
�D�[�ě�y��$&�m��N��U�OPy{�I�yV�|�q�4J�N��QXDhi|��z��;o7/����+��Ѽ�އ�����	�8��rJ��u�m��%8�r�gT)�Ħl	�XT �Jq�� Fŭ�Ɛ���\6�o޺l@ߒ��q/�J-7���F�dm��|��%L�&q�rzT��|��Hf1�0��?
�j�xI�C��x!(*���Xq�_���l@��Ѱ1�;8̎ p�l<���� <x.~\V����j��B עEm�,�2��#����X^��2�)�\���8�O�6�l��J+��AN����h�v�`~�q�Ϣ�,����	Iv�d�vVO!�D&�GM�$Ҩ�3��;yK~W��W�0,�B���׊�^�4��o���0�ʯ�շ��KWa���c���*��.묗B��C�p�T<�����W-�����;�����O�V�gj���#�Gwn� �q�'8.n�I���,�f�B�ٳ��^k�!���X&�������/a_��\��8�/������]1�
�����͏_�	��l��SO7'`��U�ވ���\�/���)��s�б�O~3�s��-&L,����~���0��SOq�3����wbr��1�����޼���q���O}��V���$��`�P�&^7��I\�w 5�lxEH_X�6v4���5#����
@k{�
���PV%8����6��Lp��~j��[�23�i�`q�Lˉ��n�"uo#BiF��񓚈e}�{�I�|K~���<a��eM���*>t�O��cu�����f���y�g^��\$�I�M���p v�Q$K⚯��a^�~�����d�ŕ!5��a��y���
T��[x���_��� -���
bq�1�}�K�쑲��h?��~�
J�&i��1�v[�媃}˰(�����9�6'�ªɓ��w}ַ��ı?���g�����╖&���lۉ#���7��NDsb�W�G݀1�h˯t�����ï_���8桫���]~����Ux�W<�Gd]~�)���q���gb���..\�e�����[~�g=+M�[���_}�Q�U�~�wn{�����g�./���2��6�W����ۨ�t'=��~`0���$����0��?xBe��u�m���܄��"~��C>�K۫k����ȳ?޷u�����{��'m`�©����0��N)7�*G�ip���˶�����N�%�f<��Z� B��3��[x����6oqi����0�7��:ڎ��^�XQ��X��,�� Nt�?3��̣��RZ����˩���m6Y{��2W���F�&�@<�+8}- ,Z�t�1�Σ�U��,t^ed�VNwL�{���$-A��o��k��}t5�
��>������^꼺�ܬ�g�{z>��1+%��e6����"I�A�T�(8Q��D|a�.#j�:n8p2�ov6 ��-�6� B!f��oՀ��.;���(Q��f|z����<k�3�f��x�8�}���-�p	:"fq�b��9�
�SS��nР�����
O><r��N;ͤ��q4��f6��r�����M���A��Ց}f� WwD���$�ú2�@,�<ħ��Cx$;^�(�Z��V4\I���U�H$:�S�/�1�	K��aD�D��W�.�Q��Ӱb>�)q�PF�o!��Q�[��Q���� s_���w��4�����]�񶨃g�{^��DO隠�Cp'}m3��M�Y<;ys���G�� ^�g�#��)���c�m��I'T9>����&͔������Y~1�d@����r��1`�~�UM:��ğ8n��m5L�t�[װ���+�$=�Fɕ��Ǚ[����=�/Mґ�G1۸�6�1�X������	:��9:~,����޻�|��k�%4s�����]5��f�����o�׼�d��__i~�{DN�gH��ӛ��Az~�y����W!��ٟ�Ys�ʣ�(�On�V�}��9�^�]���/������bB�`�5<jD.�:���f�������_n&��O�g��uV���+�GLM5s���ך��?9��#�n.�vy�.a2U�*voסwV����9>/���y�`�1����\��1l\u��}ȩJ*:�&X��?#_J�ڦ�q�c[았�ln';0�a�Q��#���}��H���t�M��MS����]:��!�@L��YPx�q���*��,0�j�9��>.h���}2����G��>{�<�H3��M��A���t���:�+=�����9i ���]A��l��0yj����.��r97��gb@/k�f�A��4�N�č�����KaI��^y�G>)�(T��|/ݒ��G�4��uWv��m�Z�ÕHQl!`q=΀ub�ý<��(<�?���U��XmNs��\�8����w�Z��	��M>+Myd�]-P���qY�&�5��)R����^t��;�n�P|�?H�E<�$�7W"����3���8__\\�ɗ8T�R`^*b@�)x�F������ �v"?��>ol�˿���x�M�P�OS��*]={�"fz��VY�PpH�]7
��~���zh�X����g��-C|�,�m�������4o��;�su��f;$.�Qr���i����|l/�P0�C�Te���|ڽ��سOrʝ}x�u���0o��]���cl�=Ʉӣ���!�9����j�~��������ܽ���is�f�~����;�uL6u=`����E�t����jT���gz����,�Xo�zx�w\8n��$4<*~Љ�#M���� �FQ$��w���n;d�Wh7�x5���8�c<�AQ�)�&H��J��N�����&](x-�u��[�EF��7ئ������3�$�϶D1A�W��a��୉P*�rES(:0w�i�m޺�ȗ|�i�8:k.�E(Ϻ,�h�1~5ݠ�#�]�Z�Ε��*(T`Ro���7���kx?er�*�$l�������?�!���oOKN?d����G�[���TnE�k������cXpu0�P��X_��|��Z�LYZB��S������X�6D��Fv6���u2��ȏ��Sp����x�t@�籡	]���x������Ȋr,��;h�^��B���B��zW�ʿ�|
��OT���V�J�}RX�Oqmd/]�XF����²�g@�fn��8�V�81sEx�@�gI�j7����>^���m�2�3�Dc����jQ��,�˿�+�����m�C�V�$��g���	h9��Tx���Q~�׿����p���N��|)(�,s_�
?q1�
����}��a���6�t�㎽9��ȍ#M���I�uO�({��/oN2�̰2�~�YL�������F���!TN�:�<��As���6�'��~��a�]]]�I�n6նTg]vюg9���LJ��x&�{)h j��»_��b&����QmOƙw�e Ѩ:-��ǽ�ȥ^���ߦ1c��)9�"����~'�E��WH3��)�͵��qT�&�����z�q�&�����yF����6��|�}���2@����g�Y��nj�$ʢ�z|��:s��{Mu���	��a�mA�:�F�����
��l�ݳpD���\�5?�lC'�k����M��`kk�Q�x>�a,`�&>b��7��iNЃfckl�\l��6�X�۸K'OD?���X���P�6�[[o%mM	�����F�>������m?�C.����K�%�l���3F��K���ߠ΁T%�f ��X�$LA=W�s��v[[��mCq}<��������ɴ0I�*OДD_Q�Fy����i��Z�OM�u�_�M-�I�����f��a:�q��x���1m9�ͳ�¯*��	���U������a�o=�52��iu�gъ�/�f�'����*}~�Z�0���a��Y�xN�7���6�=\�eV��܇�p�,�T�}Z�M�Nx=�ef�I=��㭹?����.�%.��#гB�Ȅb�=SާӃ�wXuuB�j.�=����:��羭�ͻ�ټ����_��/���r���(���X?�
�|"{iΙ���eԧ�(Gn�n
�Ʊ_��]�������_i�O�r]�^����U��X/�g?�
���`&qb�����,��_ũ���W���t?�J��(�=��j]�u����\�[�Pr����
����0<��g\�3	��B�g~+P?m �2v�0y���~עMo�v��v��9�D��a���q��x�U����e�"��i
х����~�RO���S� ��d��D8^�z�ɫ���#�6O���6�8���
�i~:�
�k�$��t%��h���
x{9y�G�� 2h\�Y��ڦ�x�
��6��z�t��Og�~{-O�B6��?:�QA9���W?����6̵��4�CS����,^���+Wi�~�u���J��<�	�����!y��=�0�P�	T�v8��m"��7h�ՂE�*ݼ}���#�w�'�9�Ma0i�, �[�  @ IDAT�3�.�<ˠ4�]
4���Q3�ҩ��&B�(�'��Z����ѵ�A�s�j @��׶޶��?�àM('�kLh�o��&��Y������܅�����?���F3�̢	g����o���k���皇/\�8Aa������B�}���͟��k.���5L�<q�>鞉X����B$�[����.�mV�1�qB/c�dk�wWꬫfC18�osrOFH��\�%�ʁ��1�:����.̏��m��I� OQ�أ,��}
;��x��F]�CR�40�FHX��m&
���([�iWy���3��_:A��v�h9a��
��:�R�~�y�Z=�7���]�o��pf(\\n��K�RyM��a�'�j����L93�5��q����9ɑT���*�]�P�v��&��e�¾���0�Zy]�6?��1���f'����xC��|��W�4�;�g81r2q���͓O>��G�\�]��D�G�-��K<�P�O��̷ka�I�B`��']xR�����4����<(�1MYGy�y�����Aͯ4����v���&� ��I�'������������gԭM[i�O�U���O7}}Wx�%��{�i]7�ߐ��@���8<�)�9��bU�N��M�|M���n��څ����Y�J��S~UGa�8�g��O�g��U� #�+����(j<y�~Ns��&������6O>�%r��쉗�e2>�*��ez��$��؇�da�U�����7W�\kV�މ��sp�=���!�����C?��ƹDt"�_+�mk��</�Ld]�W����kr����"���u~��r��_����&�'��^H�H'|�����w����az�8>�K7����?"���t󴽄�1�q�w�f*�+<��l�^�*��64^�]�^]�vL�� t}7��»N��|�X�y֯*0@�2�� ���8��8B�VS��TJ�ќ����'��,ht4�N,$�@�����4թ
63)�}������/7���~���q�7�p�����i�.�V�L���q�=�0��^�膟���	���2Z�R� S2���-<�Se�� -�A�{6�~�B�*v���ao�Ԯzg�VC��K�ؼ K���o��A�>	�M7`T�x�#۴u��2\X��-W���+W����86n�놇]u��t� �2����8�qt@\0�~[!.VU�I/b��6o?�c2�\Z*ϻ�;W���1�;�IѴ�%haV��`����*y�9�����(ë�f�e#�l��b��7�ΝZ�
7b{���o����U6!�e�W��%@��|c����a�����ؔ�Ͳ�r�oq��+��ڞ�n�r#�m�
=��󉽉0��g��7�Ąh����Ө�s�B<k�0������s2i_�l����# "����MhI�I'�U�kҪ����Y��l�a�B�O����c��5�u�09O;�/��t� ���ia����P�D<��D{Y�D^�B�[N�Th2�C�E>B�GȎҎ�)������)o��
$�g��J������Fz�i�e;��	z���iO�L6��\J�P��&R��)o�/�ď��$��	�aT�pL<�̀�'o�_qo|']�ՙ��[�BL6� );&Kdj��$÷qL���8�i�Y��|���b�����cf�z�����f䩍3N��O�I��������}�6?�vr"M�<�lG\�P+=��Es�s�T���9'҈a6�f��'�T�/݊a�\|�g���ς;
����J?_�Y�i��f}��)��+��6�<�v�����l�g|�ڸ���Fׅ�|+��G�n܊/��?��|�{���섇%��?���&�i<W�4Ѵ�{��99�;�Μ<_��>t���c;ΩzӬ�:Y��:��8\>7m���ZSr_�J�#&����3��QA�*�:|��!6V��L��p��ʒj�<�zH��`�[ֻ�Qr<󽋯~�6��ӯʩ���-g<��0yr���i)��G�x������.��)<�0��}�4���S~®��o����?�M��{��/Q�J%p�3_���©+Ⱦ�[��g��\=-�#]�,�����t�ge���[q�mŢ�~W�#��� m�cS��t{��7 �*����ei�r�ß�3��*ӄ�A�����0�jl:K�:����9@��M�?]��w�
&�5�Dy�w��8�h<��{�x!?Jl�#��K-~�g�y9����+���1Oeu5�U��G�t�uӦ&�?�(��Z�[l�i����O4�>�(��Ǹ��M4q�1Ȇ]0�w&�f�����8�>wj�7y$.��θ��5	�����+}E|������/$5ѱ�db���
���&��m�J�_T���+�<��fB� �fA-�V��Nӗ��@z���\D�M�������A��Ξ|�(Ă�%�<���WWM<�'�JYj�xՔ��-=vtS�x����JB���q����ӗ�����S<�c�t����WW�a	2���}���FS�CS�*����_E(U��V؍nҚ���s�
e��>��x�ݔ�_ij��=}������ӑ���I]�+b�iF���kWh�Fh7��ؤ���,�D����E��5�Lٶ
��oz��Ч�֊�	�4t�I��T����s�����]�`h6I<��.�co�9� ��pC+�XkL�,Nr,�ٳ���
�Fmm�8�d���ڧ�:���q?���S�4��,�����}��(U�*��:�n��++�w��i㛧��N��v���ȗ��'�uƳ��Ɵ�;8L���c�~4�~�ܙ�.��F�����|���m^{�+����r���M�t�U��:Ŧ_�c�\-0]�d���{L��P�^?��c��U�����4�O���}�,q��8m��/\�ċO�\��o���}��ú�4H<蟴��D��u��.���wa2~�����,˶5�?z��';v]�q��ݧe�w�W�F�����A��i�j���ע�Fg}l�S-e콳���
�wi_��� ̂i��~"O�Ҳ�n,c���-h����I&$������Z�
{���li�U2io)�v�"^�����'��xo��O��O�M��i�-#Nlwa4L|D޻�3N�W��t�o�.m�/>+��+��l'����8(��|�{P���n|�t���Wq"���c�*Ǩ�Wz��[�.����:U��]~F�|�;�{?y���v]B��b8�
�U<�@%R~����ـ "�:Df\E�r�]�w峪sRm��Ƅ�+z<� .�ǭ�>n��-��+�L�Wdd玲m��'���'2>������&� QI��r��Ň~U~�cA�����Z�̓�(�_[������?�Ry	{�1QS��F>�u���O� $R��W�^!�}�~�ɀ�ß~ܨ1��>��#�Γ�N���o7klLS0�vDa��><Y�g�
���*�~���y�l����~U�j��׃�wúi*�&O��T�D�*�#����QLQl�]�dW�=�R͚��N���p�{0�\���}ȆP��'�+��S����̞,�[��-^M�,��ۇ��S���	�z�Xl4��$G�
�&�&�����yly���E��ըz{�&�qݢ�bp��m~��5�p��V�u]ʛ�e�Hm<pr2�I��U�q@]NQ������Z�G �0Q�Xᤌ��8���V�v_EL~P'�|h�����KT>�@:tr��Į���j�F[z�pB}�;9��Xg�0��o[J�y|_r�:��Q��E`������[��k�j'��j)���%�,
�"L��0
{aS@5O�Jz�`��B>�ews�[�m�X=�c|�\�p>���e��t�ۗns4���O���%6�S��n��闛���bl��Hc7b���ܺ;g�or����׼�,��Ak���ɘ?8e<�h�x�>��8�;��e��"y�B��\�Mc����i�G)Q^�%x:v,�u�縚s���SO>
���W_}�y���w�}7&����h/������H�)��_g{V=�������L+��Q�8�7���^������3~�mY�k�e��y�W+�7��q�Y��/�~5�(x�Q�����ߊW��]OޗV�V�n^�/�]�ϫ�Y�kCy'(�.�K�H�P�T~�O*fl��O�z�v%��n��}�6.�J���+�����u�3Oq�Ǫ*?�^ڃ/;Q��6X:���C6CEd�3'������aB�s��@�<�)��AY��Cg8zL�G��E�f�ʨc�v��=�55I\�yr�x��������_����G�I���oiZ��WO�*M����n����M<�s�鄩�׳���~5-�몮�a�:��x�zY�9�W���We|^���p~�����
�}j~J<�F��E��E��4�+�ǰ�E���Dm�0�
������W�
˱"j%eB�1 )�e��@y�e�"@cV>��=�ر�E��ӕ�*��v��mD���
>�]x.����
�	���u�Ε�C^�<-D�k��<� ��'�n�?���a�+���=p�͊F,O%�U(6��ɖ�������e
�L�����q������[Ll��8ˇ�p���u$���{/�o<���ɧ.#�6���&&�`r&��i��μ�λ��8��r^/�.m�	�z�7�xjBu���py7�x�8��^�>��p�%(h��V;9��g��h��i:iLM�m6�	J�o�M���V��O^�~#��􏚳��?�7���r
�e./�n^�8��٧�i�?<��5��ﲹl!dc�D!��/�� ��`�U.�{
ǂnc/�)�WӿÉE�o�
-�K�b��yg��16��l�5?���9��v��c�qY�ـ���ܴ����=����|�~��|��s��~�s���Q�-p�5L�~��5O=�D�����khֽ�[�t��;���,WYlP��wp(.���� �	����q]�p�y�����tҢ���΋�P~��⡜��nxT�`.��]���t�=n/M�m�������ۡ������!��b�G�ߍC+{��7�~�ة�_z�\<�{L\pr,&���/4������?���ʣW���$�}�1a���6���������ms��Q��_N|P�pzK�g�R�)���C��l����&�x��X���K/��*�N$l�A��^~�+�y���M�ĄX�o��O�;��/�>sl*�u넧9Ͱ7�<���e&H���4r׉���rg����F9��My�K�ur�^�v2(즳��y@�� ةy�(OI7�;Q�qO��^���M��61��e��gZW(�֜ �Ŧ��O��Bv����anY�n|����>�7Nū�~[���}�_ůg���{�+lG_�S��^��(�D�d`6ѧ|Z��@�<G-ûa�y�"�]��e�aX�~�V	k��4�Ԁ��ߔ���*�N��7ƉNL2��*��đ�TA3�3�ܬ���'1g����W-X�
an�uh���v�Ryu��X�#V'�{O�s\zW9�c\娵�Y��<G๦�Y.�H��7��F�q����v������[8�|�/ڤ�[i*]��:�W;�����`��|V��̂��S�U/�^x
թ�׳��}����r���ab�?�l<F���w%%��o��oy���C���UI&��cJ0�&�]=�aH�s{u�}������؊�3RWc'�qF��+�ʁ�`6UV�S
�ʺGW0T�X�?�v�y�]�M|4+��K;�/�*o߭go�X�l;Z�Qi|V��秿n�����(��3��O푰�����a'��$Bo��z���No��F�_�j�+�]�~󧏉��I��?]	���;�ޫ�I�*
�><��R���_˰���X�RP?g;������r*N�� ��_�ʷ��tJ*���V�Ն˨ff�B���]`��� x�R+�zT�'����_k������Sg9��;4��
��әxp)��[׹��U�KO?��~�����A}0f-����~s�����'ﲗb�y��e̙X1�=����dA�������߅ �G�Gͩ�i.^Ԙ�!�c���K/5op���A��3�4'ny9�l�8α����o4�����2�9h>�ps�8���^��\��ԏӬF�/��n������Ϳ���
S��]�Y�v
^j�W�.7���dc��6�����~/����hj���t:�Ǿ�$���>��cĿ{#Bxu;l�ՙ���K�3���V���K�+� ����k�N�0��be��`����L�&I�0x������a�a�sSG������{�@j�<����'1Oc��u��&cj��9]����S���9����P��6�1�o�Lѹ���+R=�a�����7g:JoR�9�٤_�	
md�� ����:ၾ�ĥ����
'�Ҋ��ޭ��U0�7���l���e�i�wM�55���V�r���<�����L<e2���s�����?����_~�YYϾ4�{��el�13b�H����0E�Ҿ>��ƶ��)ד�gփ�j�Cp��Q6s�D�A��L:�[�y�C�Ҝ�oW*,ׁ�:�W��ʤ�jNh��$^�Q��x!��u�_O��:��~�~�0���g�[']?=��,Wq�P8l:��i�飌6����ໄs�0a0/����O?���x]X�ۇ��c�N~!�)���a�/����]��i�mh�9Q��m3�˽�nݎ�DWp��w���0&���G~R��Q��-��k�g���ϭGuW����2����G*7T	���]���aa���s�G&O�j�ni@����Qq�ʐ��g>�����U�i�gm$/0��p�V�S�B'��#�Uߪ�`T}�K�W7M���z��ྫ�}�_य़w���rI��6����O�������S�$��g���M֒@?x�[aѭ@��@��z�y��H;�\�Ce'�H�����ﭴu4BnF��j�R�[��X�s��g��3^ �'���s�K��Rh Y�).�s��фzJ7��1��ǯ%� v����^+	��>�t��$�����0`��#�i����;{n����Eĳ�R�C���H�=Bq�����%^	�Z /��4j0�|ď���t
Y1H������;�Ǹ���l0 ��PK��̈	v:��GYY�7Oq6���ؤ+�����i��0�i�qڈ�8����=6���k^�M���8�b����V��އ�q�O<��7��0�n>�v;NR��,dMn���c%pM*�#�����`�+���#�S8�muA;�V��ֹŻxs�vRHۋ�I��{��2���	��¡Pa�=h�����([����n�4��ߠI�=���EV8�������r4�~�������$mz������\���,�jV�@GeB�{��8�h?{��m��/�?���[Ax<�đ�T�	o͜�iB����}��r	;�)L�4�;ɾ����s4l���PƄj2��{(���YM��g�^�Jdd�Sk��� $
��].<t�D���Б��iG�l9�@��@����4wa`c<��@M�{�
���]�8&�ӹ�*���Mh�Qhv\AM�w��b�'9�G1Up��_�_��C��� �p���i:h��$�D"������8��#��:m��=�M9�Tm�6��U�7u����?�r��j��x��wnP�`�)�y��B�x���+��!�m�Vrb��7qϲgixz�G�D�'�?���x�d�;�ϸ�06?ٜ�x����I^�L�\=s��{D;k���qL�Ξ?�P��Eۄf8`��4��}A;�U������m^���?���F�C��.7p{z��]�'�&�IiS����v�f��,���%.���Q��<|�'��_��^y�������7�j����=?v�mp'�U;��$�|��;�����P�!�g�67�;B��A/�N����w{�7��Ɇ憞��s�ˏ�a��C[*�mSo��p�a��K�	'`:�P��^=�B7ä7iкH�£���q�(V�[%�e�����ѓ�q�5���K̫�'���F��K1=q���B��Z����W���&��o�-'~
w�E�0
?��dz���~W�51�۟4x�}f�\�8�O�������[�Q�X8	�@Z��9���r��Bu�;�$��K�8�����ω�����0�I�z���e.o6o@���8L�7�����<�P3��V4ǀ��qp��e��+�߳�:heu ��5��T~@Kީ�-��1���s65
�qd;j<�(Q��3��� r��Y�����ӛ�E_�6eu޹f#�&�Y�3��n{���������ý"�U\&�1��=�Z��H[����n����.�~�W���D��sN����r�)�~�.���v���Fä_��������9��![�j2��äyP�� ;��Ux=��~�/�ײ��DcYvv���*�x�+�z�=�w ���D�ӉP�
,���̲���m� 4�R)j����4U�A&1�;��i\�4L�n�v�\�ep�Xt�>�!��a���Wց�)��j��t>�ů	�u�L��C&d�/�w2�dF7�K���Q��I� Wtr����ТghP�#�~��!C�y�6��:!>��S�����4?��K�U���ܰ�Ч�̥K�\���y�Ye��D;�w2�cc�58�uQ�'��퓦<V}���6��<�+'N�N�ë�)J$}�|��"��Ҟi��9�y6��K��As��m&`�@J!P�0���i}c�[,o6�����'�Ep||*Oq��z��)%i��	�yL���q6t�K���hNǙ�(��C[6�y�׾�L�f���	L�V8��޳L"<�����K�?8�߅I�B��\���L 5	^�������n��o�fNs��	@�v�^�����񿄦���<i�Ʉ�8[�Ɓ�=7���_���i&('��f;bW�G��́�w�V������6#�+��b��>�����)j�=�)5z
�-���:��<�w`��=xG}�)�G��|�gя<m�=Ak�;n�>I���O{�-ڸ�Ǎ����4".�t+����������h���\x��K�K�8V۾��.i�c��W.Gz���֤џ&9����[��4���|a���;"�9W�"��<B�\K��R+��]�=5j\�*7�ϲ��$ɋ�Y���H0¿O�5&�+��\��Y��h.�IYrK�IVc4�RA�����?߼��k!pO�H��r�C�9x9y� ��0T{Ex����/�q�AU���W{W>�]}W��b�A��G������3�����|�o�W�Y:�^Ӫ�K<S����?Jj��:T�Ȥç�6��tm����B��(헚0oz�2Mo�Ug��QPv��7�o��[V�-8�[���<u�����7��^z�G�b�g��^��I����x����q՞��suкG]Y%r���|�+_	��x�#[q��������ӲB��U��%p��-���@U=m6��{�˔���9�zy�!�`�����5���%�2����/,��K:�g=��ŷ��+2]7��|M�Ϯ�p��a�����g7m�fz�8�����mP�Q�*�ϟ��P�&=�x��q,��f�La9o�ͼ:�^�}&�/��2e
�$P	H��0�$�b�_u�"�|:H��@�?��yyjE:�4�Y�,:;��ΐ��"��K�p2:�I+����og�ߎ+� U���e�D��ߋ�\�^�c��TfZ����'����i��o���,�_'
:�+�Ǡ��i��2_5�î��_�G������c@pf�ω��1Uh��Q�GҴ�Q/��I��Tx|�SO<g�o�e����hS�v�l���o4�<�D���'�$�Ż��p�����8ڣ��A�Ba�aS��<_����{������q"�-ݦ�o��
,᠝�9��?5�_:�1W�r�Js��C!īE[����&��
����M.A��w�k�/~�s�ݤ9���iJ78��Ϳ����ʤ��<I	,d�߻I�M�L��7�ߙb*��J��s1����]N#�ZFdQ��j�g�1`3��hf�u�_��I�������c�b��4ǶM�iPgˤ�
����CQ��VŰ�=��1���Ӝ>4}��[h��_�&Sj�=R9c4��e�ߓ�ą4�<��{�������_{����G���J��k�V��?'�)�zc�qķO7Q��^�')��ֽ~���i������ef���WCj����|�:5���k'
�
�ބ���Ӎp�O�E>��"��nM�S(�;���[��t�������?
Ws�cBڅw�땽�-�zxɢ�m�}� .b��$@S3�FX0I���{���sg'7�o��P�W��l�-�VŮ�>�o�p���c��o;�������ͷ���l^��ˁ#���m]�����g�: ƘlP��8r������ɧG�W��/Xv���@q�_�ux��W�4e��ч�M��Ӟ�pB%�]]��ێ5v��0�]��WUf�Ix�+�,y_x��~�᪄tp������[ͷ���k�<r�IM���G��m=t����g[���cI�)��.`mۦ�Y~>�#~Z�S�t��)x�o�pS��O�G�&p����js��cy�,ҴyV9����<U��_��m$�O�W�o]���g�8�~�� ((���xJ���Y?>�b��v%	}ƕ�1&$*�vX�l�jE�iF8`a��zw�&��!LQ���N��g¯<�zV�iu&+���O���������3N7}�[������;���??�m�D�m;]����?ۊ���_���m�.Tf�'��~U�U�EVFE狊Pd�V0�LB{0L����LdOH�E����u��m4�qQ bx��"p�b���ӏ��b�^F��\� �fMx�?���{����L6���3��r�"�p
"���컗:)H{+����˲�9�F�io?��5��vd�p?����Y��av���m���Ε8jB��L4,����\B��:a��9io�i��s�Ц?�|��q��;+�O^�q��o<�<�I-nl}������\�`F�;���J�I�x��+¬xZv�矢���v�t�����Sc���
�]��\��Ɗ_��oi�ʐ���|��{��c�jl��X_mvi��I6�"�y�Ú&��||�Nsgu#4���,b���������o��.B�ܔg�#�21�������L2�9�0�pB;�K
Пf[n��AM0������+Ҙ�u�F ��]���
x�a�w6�ӻ��ғ����П����?����U�g����u�G^�[�'W�~��p�6�n2y1�v�W�U�����ʮ�B� H�Nj�`�~�qª7xP�<	��!�!�
�#��u6?�����ǓZ�uֿ���4��	D�y�Dv�/���x��	���GF������G��X%� |u���^ >�Y���[�f��Q��&;q��y���=(�'�(�e��m��Ʉa���D�:�Fz�ɿw�(�-�����l�W���`��[��`Esp�+��ɂ8�$o���[ON����_��ƅ/����ފ���+_�O�����������|�.�����~۲�`O� Ao�.�<a^T7��:����h����3^�	���J_~�q�������62���]��&O�IG���ě�ں��>��4}�ey���QO�T>�e>=�)��ǿ�������M�)��8��C�u���nԱ��+>���0
ͤm��w���!?�6U�K����J��ů5o��F�!��/'������\�d�ū��U!'�/_����0'��w����yW�70I�4���ܘ���!潟^ǜ�~䱱�o�phY*,���a�>c�{!���؄��ac<�0�r�:�e}�Ϻ��~ґ���҇q�/$߲�ҚO�&ϯ�����o�Q�6��YF�L7HS�����t����%~�t�:T��@�^>�۪(�MJ���V�W7�n�_�{y��㐓�{|��I�����-$�S8	mG�WF��퉐`#!��W57jye�aw2����*��ͦm��U^M�9�<]��AK&,Ӡ+�9�>��e�V��HllĎ]|���p?���'��S��9��`ƖB�E��K!t*8���N&%�1����lS���#���I�Y����Q�j�՘]�r3o��RN�ȫ�e
��X/�ϕ�;��j���_�hȥ�-V.�9*�U�k׮6�<v�y�k��|�C��9�¾π��-bϙ�(n[�	���TA_���U[�^$�WꛌOF�qG~��l��g��ğ��~��I����}{�y�W�ϱ����Μ|��4�n�s2v��
�E�G�<�)/1`��h���,��j���\z&���Te���k1 �����~�I�wïB�����Mʱ���������e��#�.��� �88���+j�i��V�O:�4/l��+�FAE:r/Q7�SF'��t�Ħ]�V��I�~��(���Y�ِ��`k���؀l��yll��ֈ�~�G�<XϨx����6P>;��ͼ��G���u�<'0Ҽ�ߦ�TA�|�1q˶�}	��i��n���!�����.~rls���v���㹙�8	�	�yS��UG:aM�C{/����囯uȶH�u��	��0i5x*�����fm�qm�����C&l���\э�i�'nl�#�¬�<����N�	�B�{*K�1{8�@Mcb%^9�,h���lca�>�d��D��y�o�����h^DI�����#�!��]Y�b���ϺZGW8u�w��'�����*��N�_�q|7�~A3�M�s&�A���IEќ+v��R!~���E���O����<˰M5�i��'>�^>�'�7n<i'vNn�L�~�"/Z1G$���S�7�k)��e�Ҧ+\E�j�Ƿp<ȹ�Qgx�(����8���
�m��d�6w;��˙��^����(�l�Nږv�O^~����7���k�g��m�-��� �[7Wh��T���%.�s��>)-;���1�%ar(�I����#�	ƚ��׺�Oc�%Nե�G"��=�����_������2a�a��C(��kX�n^�_ê��[����w|��2t�_��Bx.��N�{߻?:���7�nL���U�W���tP^�г:l1����մ|�,��Ui"N�>�����pC�Q����o����1���+��pj2��*�Z�x�͂�AT'C�&s�����'�a,�� ,���^�3�M�vD�UWWN�ͺ�Oܹ"�9�(j�}����\h�ꔜ0{B w2F)]��?�����Æ��o���Sy\
����͟'�a��!§�{��£gl�`-GF��A��ͣO=���_{�y��Kͭ7�^�s|��f0{��=���[lf��!�|1X�_8p�u����}O:�xƩ��t��U=�/s���«������I_YF���h2��.���w���o�7��\�t��sk.��u@�M �p��:���H�	K��#��&Cp%m�r��&8�궱�5��e66�@�,Ǯ��b����e�.:[	�X�]-����yP(@���E_P������x������$с�L2čZk�9.��V�{��Xiv���q�����f.�s�`����F�t��|7��i�G�������D�G���b��dO�:�-�^$�j�Bi�&\�{P����<&QӜ�d}˄C��9��߲bb�N�l����1'6R��dO8��c��׹y�h籫clv�e�2��&C�_�O9���o5��\^fp ����Xa���g�ӑw��i,Sۆ��)J������KE�)<�V������K���0'0�9Q0M�ds���`�r�1�Q�!��?��;iR�C#��ЅEO�2_�	,#�f�ܑw@̚)�{oݺ�|���o���盗^}��1�tO��t�e[������4��w�tI+>��?�W\��Mk��ԍk�J�Stb<�:�¶�[��O�lC�u�yB��rd�lcaQ ��3�z�Y?�|/8����dP:���~z=�J'��Ε2��楫�|�K���oeР�W	���e��
'����]<�&�7˯V����Y^�޼�������?���d�B/>�z����X-4?q���w�#�� ���C�s�q.�Ұ+����ǟ4�+(2Xo��k2܉��z��C;���/܅7L������p\�fbO���7#m�����8nUi��~��g���+��$n����;ê���p�*_<Vߕo�R��������L!�^}������0P���������Ji�h�~�"�����N�}�����ID��L�Uᆥ߀ ��3�)YE�� �+��H�35%�{��������$��r��a��Ox���(��<�&�K��F;�G���m����+�D�- ,$�-���@ffgY��>����|l����ֿ��X��M�HJ.���{�����'
0C�[5��d�A�)�=<�ģ&�L[m�>���E��m���a�[|:G('1���O�"�-�����N͎7O<��&��z�Z�2��Z��+�uM�7��{J��~�3��%�z�hmC�G�m7�l�WP� RKi���@]�3��iR�S��3����o��o�z���=�~xuKWj��d-�0Шiew^�`�u
\*�Nc�cYnX�d�V�ps�B���q�C��0-A����$�����[l w��pjVvt�>N��ހ�B[j��{�i��1�kr��5q��ı���X�I�U�8�_Ls8�s��.�;х~1��;�C'ʓ�������y���X�Ci�wq -�n�7��R��NA}
�.�dӷpe�����R#�tW#��愝�r�ǰǊ�}����'�9i'������4-����*��n6j��Ӵ��0�-H���n�1��=���f��'(�-qX{�*4u�n&����=6��q��\K���v1;�nf���w���B�7>�ث������]���m�4�	�eXW��M�ڮ]�8�3�՞�#���e:�e�v�N*~�AN(�d2q�Iψ&}���DͶ��MB�ru�f32@�m	M��'I>}�Yv����~�Ն�CeS�ʓ�66�6'���y��ex�%����X�u��>��C�a����	�a!�J3�+om��[��&<Q���O~�i]�����C�0����U����������J��4�hݏ�l��t�e�9&:�w��w��ֲ}�i�-�8�講?��Q/⛇�ؗ���4Nh}7�2��>��À_������0+�L(��q�[E�͛7��N��P���W�������96��t��Or������53;o�$6��wE��c%��|>�J�#����x�'	ʃC<io\�c�<R�p�p��s�ޣ���FWO����g�<�q�\�T�	�n�����g�o��麂��4���w��S ���p�n�_��bxN˯h�r.��V
I
*�~�: ��_�8����wiZb��}�L+Э����+��%����͵�u��  ��3�'�eY2;X0,2�\�r��BZaƸ!�0<ӝ�,���|��v����8��[�р�qT�r��i�t�8��Ǘ=T}G���	�B؝��䧦N6�}�kͷ��-M0̓���m��$�̷�_�P�cC�wr�Wn�1b9�U��Zkj0>Ƅ�r�a��0GPD�I��9��}�sh]�p?��B�En2ݯ}�כ�~�1��{��-6.3`�#�<������d�\uզ��~7����~� �qM���4E�=�6˨tN�����l)�9/��U�,5K�����W^l�]���Q����3�xs����q\��p��K;�#Ī��S��1:.��S��fJ�=�]�n����D=�x����܋����;9 �~���D�z��5���{�$�#j��v���w�X�P�	B�A�u*ܾ�b��f�&�A��&�!��',
�^����(�Ch���\����#i�]A�>�P�iu�{@">��S����%�6nTW�lP���������  @ IDATʋ���p��-Y7�#�*���L�Ɋ�ƉMВ+AN����Ba�G'B҉{L"  @߿�ԏ�鉩_<�N��U擂�{p�GF]�.��Ŵ�쪍e���B7	9L �f;�{۴�ܥl˒����U�UЏsb[�D�i��%.�����Vx�q���w�|�n��J	�E�����D��q��͍mB��^A��ӟ�:������8��#ܖ�u����k�/T����~����l��[W����T�F'����(�7�{y�a�x��X�S��#NZ׭�Q��[W��G|��6R5�R��ֻ�. :�^�!}��a�O���p�V�J,��t�%�u�5�x�����O�o�� 3�F�|����D�<��1��l�x�\OMސ�r�N��[�3�����e��9� ^뺻�*�0�pO��<�g�]�|��)���q.c��u�}Mϓ��9У�u<?��F�4��?��}�H��➄Q�©p��;.��G���-<ū��Z�n}�����L�q�l�2�e�_��^N��O�
/��6̼��+?��u�)�/�??�m��<�����H� �&L�A�N���;�}\Of/q&�ޟ�p@,���
��)@����p\BuO�����kM;��G�0���lt8�U� :�Xj��6$��>�E0=MG��G�r�Ļ�.�:3v4��-�x�u�-����ɹ��דc���wP�SC�Z�	NW�bBIK�#��� ��pF���'�Q�y�7n�D�&d��Kj%j���5pĎz4P
4 >\Cc8���G����?/?�t!8����x�s?�m���Du�da�v��6}���<��������'Q˄��I;�m��T2c�0GB�f�,��w�'��:�&#Ǵ�K����X�r���̑�<���h�	3�zf�Q+�
x����6j5�D� ��O?(�6��w�Kb\�R��n �O�_z
�C=4�G�����{/��.�䮭6�����OC����!4c���!Ӻ�o$��g�e���hݸ�в�0G��AE-[�@)�)�T>վ�Ai�M�S���YexY��w����C�¯��_o���n'��]��0A�^�gf�wO$r�rj�h�>��)�z�È_^���(3λ�>��I��A}��&qŃ�:��7��|�6�Om|�)��f��Q�.�F���?�7�Wӭ���]a]aZ|�m��������)t�����`�M݁��gyc�GxF)��i����2��]?�q���~��]���ۼ��Э?�l�}ї���P���UL4�)�d�0qc�i���.�x��7��`6�bnc>2I9ެ-o􀌺W���������i���� �q�����������uw���w�m�̲Ow���;����+��C�G�c&��}e�=f�3l�{H�����#�9���m��бx��X�c��"�ω�ξ&��1�#W|z�u�d���vމ�����&I�ö4_����x��A��?�m�*�1�|��5�L�&]��p�Ӻ�d�,�	��8�����;�W}���_~;�ܑy�7A��&8��O�W��sv����_|��|�U��w���ip�L1��J�fi��y���)�
�}&�{\����v�9Ey��ũ{�s�	��6{�T&���P� ��l��Տ����S�8��1�v�4���lM���/OO�I���y�JfS��ikYFҌ�I~�|�K�d�V{�_qė�Vѐa9>��ƫ|��b�_�/�q�m��k���LB�a���F�������[X�q��]��]�����H@��<*m=�Wy|&~�ۀ !@a���z��M㒭�
oI�h
�Kdʜ�S��A�wY!�AH>uDGu�Wv���=.�J�y���xׅ�Ij��T�#0?�v�dN�A��T:����BXe�b~�W�>��S��Ѹ�<h�Iͯ��ө-��ꌯ3�̣H� ��5�+'U��j_���m��,�j���6ݛ?e2waOF��,:���^�[�.�yy�����/��|Ȳ��d8ۘ�8�7ʗ�Z��|�x_��2��G���g������L3X=3�e:�)t�{�QЃG�����x:��X�rX%��"#/��d��٘�1��i}m�bAPv��ʺ�ld���O��N����{2�p��Z������ll����<p^�S��t���g���_��B�N!%���-�[��r�Q���t
�N���	�8B��8i���/`Ww�;ﾰ~Y��>�td��~m;׷ez!�������Ar��`��[|*�"�����'Fz�����X�9q6����'��q��1.��)L5����s�E0Vx���q�t�k��V:�4��1L緮`�{�ь�������]����~���F�_��T�U��}���(?V�r%��Y���@���c¹O[���V��^�lT<�i-�x(z�]]s�B�����x$�u6ۧ}�Z�
�vM�oL]�q��7hK��2<�G��U�zV���ڥ��wd'm���'���$ٺ�Fe�G�nm�[|{"[7=���3�I���]'v���\i�j���*�*���mh���j��P��Hg�s�u�EZ�kdD���w}GZ�|F�۶$׊�~��6�e�:˟R�SZ��h�d^��ŷ�#|�ϳ�=�M��%�4Uy�4� Q��N��"�q<������K;���WN^�B84	vE^��$A�U۸}�f(q4崏����Q�ϓ��{�. 6ࢭc|!�������s�X������:��Og}�W�*����i��~����~��I7n�i�J�v�����J��U>����c��S��?ۤ��^�Vm����Pt#v�������� nG��)XUX12;��9���t�����X$3i��`�@P���D^:?�::���������i�!C�ώ.��0��V�E\MUt;N&`�k+��;�ܹ���n�7�l��:��cčN\��'�ᴅ�qx�g��7���w���<���� T�2}��ǹ��qt
8:�%�މ	��>�y�����1(Qps�͝o��N��{���
�ў0R��9����!��ɛ��t�͙��n?���{o�L�iĵGu��1��xOx-?�Z#�,���G��|,Ʃ���4)-���tM�db�"P�i*C���D��h��@��Cm�{�;��@s���M���D��]�|`F��8�Q��4"G��:��W�����[�m���;��B�ZH��tD�Q��F޴�ȓg7W���?�a/�Z<�_�����<J����2��ᙌ��W'�g\5�Q�?����B�elj���LN8�6���l�1�a�o��S��ɔ;҇)Z�&'����q[l����2���$5oi|����?�+��7�����r��꧿~D�'T�O��\>��a�Tʤ ^<dO��N��/��lۤWJ���jU𙿧o�7
�y�1�p���4���	����j?��_�`��:HcZ�EQN+�~��[��Oxr���5:: ��ػ��͎�>�s �@� �9�`�Hъ#{��<Kw����5s��H�A2M�2�(.Q"�D��� :���v��<�_4(��}�S�T�ڵk׮�]�l�>�Ol�V ����.��S�Q�;<�-�ˊ���6風ZB�*�e�7F=
��X��(�L˦25���LGB�̠8�>��vgV�"��e���2�<V8��yn�.3��5Ǩ��[�6=�S��� ?���s�g������C��9��/\�����74�~1ex�e���{�`.}#�\� |v4�α��#�GGFgH[B�t0Фݾ���g'J�nf��̒��?<�N�MG�6I�m`�t��:ʣѮ��n��\珰�6��צ�gg��0����%����f:\�q�P�ٵ�����G��@�~��[�7���Z����U�"�Z�C�H8��ҭ\ȭ�>�nB�_ES4;����~J����S�[���P2�O�P�lPn��r�¯r1�5�6��ɉ1��7zZ��$T8*�AS�33
�G�L9K��%�N�	mg�[��Y�+
�]w�V��Z�p4낫��=�|�����yTP�K�oF��k<�y:�8�{��un�N6<;g%���on��P�4&�+*����q�����OE*>���?��~��i\����h�)�gj��ln6
��[n��.�L��b�J�W�k�iV��T�#?��N����HǠ߹7_��[���aVD����Z�+�&����ʇt�;^'�0�:�úc����
T���&s��g��j�"�i�l��7f�͕w�T������C2_y����L�M�ﴋc:�V$�qi
n��x//x�gx�-�w��۶�(�Y�ntF#&|��sg-=�T�N�O��9�h�UF���8�ְ5mh7����ޙrϴ��	�rR�rn���R���qv>�AJ)���s��ʟ�~Mc����{����<�>�s��z�.��n����K)�?��3Yf$"]q��|�o�iN�W�Y;�=9�z����������鱡\}�_�Sy�4ZRE���AVF�N���/�i�*�<ݞ%��/�C�Z����6%.3��y�D-h��iނ��L�s�岾���w� �`�\��m���Yvvfd��fV���t:̎r�������:Sq�i�'�`��7�g�O��ҷL�w�`�G~,��+�?���hO���r6��.u?�����-cE����Qj���5x��J�l���h./�*l����`J���A�g�{<r�������*ic�˝8G����"��9B;��ME�:�O�r:�������n�&K��o���[�_<�h���e�T�C[�����)d�^�3�><CO�y���}��u�Y�!�ì�[������;��oi��I{��6��̇ρe^�1YU�t�$G�:?e�ƬXז�PFq���o���8kM=��!�j TV#9�/�:�SayZ��� R��[�mM�8� �/bZ4����p�#�5��)��X��x���Q����MyHM���`���S�4I�ߝ;-���sG.�ʭ��8��pn�6
��M�4.T�T|Ec�,�j�]K��w�g7��ڠkGh�ʝ2�y��I)x+>�?��l!�K*��>^r�Ӂj��Y/�RWt�t�,��_�E�=Ҥt�/����fZlD��Ԛu��$���W�^i��s�*�ƭ3!.�8tLl�˴|��&�X��*�������YS����̰�8')���(�SY
�ne���y����O���Y���3�d��G���i�R��'x�[�ʢ�\�K*ɿ���tz��	��I���qx��q�QT��?��f�-�s�;�h���\�P�㧁F+���a�?�p�GW����K���K�`�)�o�5��V��ϐŦ÷2�0e�n��o�vk��ͮ{H ��%�N9�_h'�ֆ��ntK����T<z�`s꫆��<mt)����4|�Go�-��A�Fg�A����ȡs_�fR���dnN��8��*�o�j^y!7U��,�����v�XV�N[���)!�߆i�1����C�2l�'}�<%_�b|3heVq���0����ڟ����e�C+x���i�Ϟ]�Յ�:R�Tȣ���8u(Yx��l���_�g��t�q����%)�x�(�YiJ2;�`����m���x��}S���D����3��
�:���q�+�ć��ձh ���4�biGr8�M�w�f��\����B^����.Fu�,�u���oU���9%��g�+t�<1�Z��J=q𧳇�dg���t�#���k��9�q�p���i�C�IN6�`��_0K��m7�6r���S4��)�Љ��%>�n��{?`�i:�Q��+���-����%na>2�=�r�Sߝ��۔�a�����Z���7f�����f_¥�0�4���`��ß@K�B"��Ѝ�}�H��</.�	OaϏoZؼ3��Ζ_:w�j9q�Ȏ@�e�Ե��ӘF@T('22a�De��2����<��l1��:9��bs:ȍ���siM�
��з�6�I'^0g}�G�M�J��l0
� ���G
�`0�_�-ڽ[~�~��F�i�����d�p�c1��k{*��x�p+�C_)񐟞ws����l�ֻYv�`.ʝxn�L��NvIX��37d3����pRJ�NQ�>5M?����+����aȎ�(��)��H��H��=������G�0�J�����G3m���;����kh���Vtt�}�G3Z�&�v��ٜ
��PT8Fؑ��yzt��~([���:��x|3�� ���4�g3�_?�f���S����Q��:.���,�w��c�ˮ�(�R9ym&�GU�D�VI��K/Y-1��n.��#���t{?�X�9}��~_�1����3���a�h��\�˚o�������v�AF܄�����_Is�3��J�fJ�l�^����s9b��N[���K��;J�<�89J��?�����sK)��կN��}O���#��]-/<��!n�O^v��H�N�8+���.N3Mw�U��G}�T4�0��.c6��JV�u��4.�t����8f��O3+_-�MZ���L=�z(�p5����ƨ?��c�����^�Qo�˖��=+�-hm�`��=F�x��n<��/nf���)�o�a�fǀ���p:���m���n�}��c���M�/�ζ��txv�M�8�0d�iju��,_y�D7��>����@���o�h����E{ʒgi�K:ᵼ��������R�}&��x\������pt,�[�]w�pcj���U˫����NO���i���ݚ�J���#�7f����g~|7>n��<�Fb��o�������5í� �Lr}!e����ui�Wl�}���?"�1
�ʋ�p�.!�z^�,�ˇ���#|�)F���ٮ�K`}W1Y���\�(��35$#�n&UqS&4�*�n����օ���ڎe��H��o���OL���Z��7R��E��G�E\p7���VY��*��5����y�V7��U	�	���e���u�e�С����J!sD�,�[9�������殈W3�>�ʋdC����N	��n����t.#KɅJ?#A�z��V��vܙ�O�i~H|f��'�=8qZ�Ĕ�̨��༬��:q����̧s����5�]z�?��Q�XD��l��p�X�WOO_i��S?��y�(��+"4���%x�4%��x�g�{RW3l���a��
Y1-/���!F�#�	#��=C?~n�/i�x�y���7���i�}-)�-�'r��5�A����>������o�3=���ӓ��|z�*�o*V2�iC;������z����}�����<]}��������G�~��! d�^�J[p��q!�ۍ<yq����uc�i�7F<�,��P0�0F����Ĩs,]Y�5�3�7s]�����"��R�b_O�T�,~�;��i�희0�J��fȗ:V�"?�/\�(�����=GNk��;��W]��Y7U~n�qI���ٗ���<[a�2�[a�Qglk��Q���9�u��L�|f�P�B����蠰��;�v�9!V��&p�`[�p�.�7��۟���$��_ܴQ�������8��xg�k�Q��3{�˛�A�s�ǎ(���-��Fd���tɷ!ǃ魦p���=�+�ntxo�z{j�e��K��������3~9K��cJ~���cVZ��z+��}>f�T�M~�y����� ��r�~�O:�����;!�f,,�t*�;�`�&2����"\�A�ެ}�ߩ��qm�g۩,G�(����Sn�6��)J����-����6����W�������Y�v��dP4ڭ��1��Kޘ��ዶ�f3K���xZ���'��0��f��B��χ΁Ώ��u��GV�sv��y��|- ���p�RI� �H�*.�KZ*||�-��8�n�+w��+S8�8����w��Y�Og�át ^;�FwG�s�0wt:ؔp�;�З�����f9�ш�����L�=����+k�͒(#���R��[�#�F�4�a����M�X�h��pp(��qI���,Gع��(�0�>�ѯ���5ҕt0p���W_�����R�`�N�Ca�*o��]q���2�=t/iWA�L�8��È�8RqdT�xO�iOP�t�p�ϪzQz2yw&��ˉ]L��gN��Yr�[�Q�J��f��F<�q4��~Ϟ��6�s��%#��(��ۖ=2��h_~�%��.�.Ʌ��w���=��@�J#3NA���;�g׷�t�|	��#p�J^gw��vz��Ԇb�ҷ�'�\nd��j)F��w.�~�ن[����K\�{��Q�l}�ꫦO|�ӟ��Ow�Z��#�C��}��G�7^+
Q6L���r��b��.+��vV�#s��D�ʚ����i�����LOd�����Y0�)���H�8v��?p�8�-GD3W��4N>y��i��X��s��Â�t(�q�����m��V����ύ����w_(����r����q�#�NAb�\������xz���d\��5
!�⠠%��e/�OZ�;�`���3|�/�8���r�y�gw�40��㓟�nN��λ>6�責K?>=��ӳ/�X(�^|I�0w��>3���kK��l����FiC���g����J�<z�	�U��c�m��X���r+�0hj>v�*E1�L��o��Q��pӉGWt��A��[yS���H$�NR�����P�|��cٝC�Σ���^7� �����ݼ���������}Վ�]}�����"�"��������Y��C�7�p��ܙ���.��@������w�05�0�+F6��
i��N��ŉY�Nœ�jf:x��sL���k�D�2u�Dڵ�aΤ|���~t�f��ߖ61��h-��3����"-#T]�HO(�C!.r����:�:^nſ�ɠIW�
ϰO��,ˊ��~���hh���O����~���0�psXM�����9��x�<��de��9-����U<�YEF��+��j#�J9����8�QH"���on� �B&�ڀ���]Е��gr�A�x(�t�k]^��(d9q$#gz��>픞�7%��K����V$L�a����H�q.Sj���02mf�6��Spdf"�Ŷ<�B[�/�W*��FzS�QU�pe�F�C��E�x�.���� ����'R�L���� ���ٟ�"cTn��F����xk
�5��ٕQ���Ѐ��B�tK�� �v�f�m5C�K�r�����sny�����w�]n8��s{�0EA+L�.ҙY���;8����KGh�,�����	_�G�<6��/+�*~4�̑����l�m��oy%ϲi������S����������)��Xp%�[i� Pŷ��oIy��ڤW��m�ţ�"�G{$k�#�|�tՕW���u���/�\�������]ՙ������]uMF�����I!Y�t&w������q��Ѻ�l6��wRWV�)/nT�}�gk��訁7;�9:�;�2U�rd�ٰ�:���RL����pn�A9�-�"SZ_ �Юȋ�Ю�����{
e�})7FM���[o������ӽ��=�Mp"��m��Ow�{���+��<�eh�����3�5r��]���ש�(e�艣��y(�܎=}q����K.ݓ٣kkώ�Gu %jsiI�9�7o�i���o�5�֊�4�6���L�G�r�Cg"��ˀ���3�9���'{�>����o���s�����k�����,�߮��̼8ޝ �J��L�����'�F��dbS"'�A�b.%MY&y�:G�N�yx�)�n�'o����X:B>���IiU\���2���VY=��Fyv(��_��|�`n5~-~��'��:Po�����o�Xw.M�(94�^*�!o�2�JGܤ�&{i���y&��d�b�J��oK݅o�輼�lN��U�_>��QO����:�ut-!a��w ��ӡ*9JX?*?���^�_@{�HW}GF�oɀB������K����BY��z�w崬���qx/��&t6�ui:ea`-~:3���Eq�r�u�O�f�4���	ٲ0��:�5��Ag�"��)>ŭ��0^d�ҕ���3�QO5�uV*o��{C hL��@�5#�t�Z�;T��}V��L'�Yλ<O~"k`Գ��H�l�r�f�0�#���ȿӡO��Y���v�1�JU?X�5�ة%� i�O�&�8�Ņ��Ҷ����!R[�'��޸�	��Ot]g���*��41��~���x��h�t.�<�ۑ��x�}M�� �
?�?�ߝw�&|��f���b+���A�[.�C�iT��pN��8�ia�/��^5�K�C��nv~U9�T�<������aۧ$�#�e{Z8 �{�t@v@+���7}�����ǔha�������^Қ�0g�0JPuN�yD/�U���>:h��3B>���)p�a��0��D3*��6��F�C[i�����/d6��V���s���h|;m�G~�|�7x<��wە���[U��V>x:�3��*��[�ϯ2��q0+Z�"�cԤ��ƶ�0�w	�q7�����k,�OsQ�ڍO�c�<��"9�� ?���������[r>���<�9}��?���ÿ�b�v*p�]2�~ǭ�7���Y�s���|z��g��^{-����Q��P ��Rb�0h�ش�5J���������'l�{K��/ݭd��O��V����r�^f�i'�VrP��{�	�4���@���__��tx�E!���y񅗧�_xi:q�X���{+��A�o����4�;ҡ�fΉ�3r��˦���_t������V�J��݉`���_n����~R�
��ͬߖw�'5�[���
K
80�|�͕.#�7�pC�e۶��9{?����I.x g��\'�Y>��y�>��S�(*���ң�[�����DN���?9���ɀ�%Y��|���}1�/���:�ኤM�-)���Ug�h��ӄ���W�-z�t�С�'�2��a�ǟ�U��::Q8(ݕ��.T:J�"
��ÿ���t��%=����D��D��9�~F�#��5�~o�vGw�7L��үÁAg�)�<hd�y��ܥ��w���p��Ϭ�0�w.|~�љ���O�%��!�M�-ݛ�ۏ��aX��ni{��7=ͳ���ۯ�,q�)��Ͻt,��=��x����w|�.|���	�c�t:��'�0ޗf�05`���$5Ug����5]¡�����'_��N9^�j"�4���C�CQ��B�(k�|#;-��z��`3��.��ÎC���������G�w� ��q�%�;-3a-��C��3���荑��|�oM�8� DtӐ�A[��[h�k]�2��ϣP}!%���1k!=�?��5�u��ӡ��X�B�K����z��Ay�I�����.�����l�/���<fG�W�Ќ`�!0n��,�t[�d���-W��к���woX'����x*����.|h(��RL����&��1�>�e��;��wf�;:=��='4�0�2ulh�ҜD����9��Od�7�L�mTK��#ӣ�>�5�Fi�Z�T��F����,o��:���S�Μz��<e��f�;��q��� 3N;K!�	�ŉّu��Yy>��J�cT��`m�|��m��Oz��ş�jy���
����©��ߝ ��ET�e�)�%�C���n~�"W*��Y�|�\�O�4?�󧳆��tzg������i�xiF��&FJ��yv������x�����@�n<#~fy^z���.��A?��?r�]����ne���o�3�*\�	4�1���0�o��2�t椥0�j��� 7�K�)�v�k���ع��}Q�o�������dF�QN�����_��[Ι:L�d���;n�N�8�wy��'�Q~����:���t�{�,%{%4�N�C��dsϥOn��:M:�d����G'#�4{j�8ߡ>���n���¡�
�gF\�cm�^���!�u�y6�61�.Y��=V��U'�����)E,����io|��f�F�w�f�-�r���KO�Y�৙��Q�N����r����G�%]�lz�ۈpp��?�n���#�N��6`��r~�۟-��f]��7X�����7wl�������fگmn�v�sg��x}wXv V�w����5vሌڻ!h��ȑ
4��;�¯�>�Eoa��]�7S�)e�l8���<�`Uu��)���}_��#3]gI�w�]~���N�wx�Sn�>�/q�����ǁ���������1��B&���F �C�F�=�Z���a.���֛l��xV������h�P�.Z#�)B#z�;UL��KB8ډ�p�9�sAo{&|�I�H]3���A�1�#��6����'ȷ�{�R�I��aX."�ĭ R���Y�J����m7xw~qS��7`=�vc��S�8�'�l�ޒ�/#Z�l{���?G�3\ֿ_�֎�0���`C����G6J�H80�Ƌn8�˰�y<`GcM��i<����f,yH�_�Zj�j�ҳ���%���x�ɥ����[���+�K�5�ϖFaɃ��k���F�8PK(F�_LO<�T�������M�dñ�W�۟ͮ�ax�WJ�{��k�T:3��)�N�i^kH�y�g�׳\��	��7�|�o߾Rl���/-�^{m)��}��PHͲP����;kiE����g����_ܧ?�����?>}�φ��2���ĳT�ݗ�~�%C>���L�������l�����?�a������k���{k����e��[ӏ��?�r�wq��VY&���~-g��R�X���r����+]j)M�n��ޕI��_n���^�c6z�p<ǲ�(���@#:Ţ^i��opW�2,?pM7qߔ����??}������Fx�&w2%����ߙ~�ӟf����{�t��?��?K>�_���;oM�>�l� Y���ji�С�ǟ=T��_z�JY�X�a���{�n��Κu!#���I�q�Ȼ��c�j|��r>�+}�@�l2�� ���$�yu"|m��C��t���u�}�7n�kJ�5\��\��w�,"�������Ӹ�m���;����n�Hwr#?K��>Z�ğ����i���g﷐|�A��9����im��PHf<�3���U��Ҹ;{������1�^�*��w�uX6�n�r������7>{�{��Vq&�%|����+��$]�z?G�f�37����Cg�� O�E��w�0:*H��>dk���,o�m�'�թX�S'���K�C��� ���遳�bo4+��_�n֩������c,��~~K,�Ȼz��4bV�ި/���A�ԅ��#DܗFD��K���QM��p�h��+fԣ�\�P���;�D�0�"�D���9�%� d�jĹ恰�Զ��`�����I�֔6��,GxҡP 4X��XolM牌�ԥB�w])	�p�yo�;Wf`(�'��<����E��w��n��;>6<��>*�|m���ll^S�X�ȯ�7���[��{��/�X�/*�K����M��#�}
FxF�!G���>�K3�/�V88Z�[32֚��L���J�X/-=��#~
�5�v�pL��Q�n�n���E�����>~��`?���K��{J�j��r��w����>T���7��/<��Z6���}���K�eMF�������<thGm�J���|�C�F�Q�6 �x��g�/7�a�ʗ�<�s��թ����H��B�S���^�Gsr�_��_եe�M�_��Wj�2CV����d��������� ��4}�k_����'�<�Wd��d�cO,xuz�������>}��N�G�����t�:^tX��t�?�C�w��urz�'���P��=-f2�(�W�[f�\�t�,:[.��=�u|�za��������[�>����؈��fiR�s�����O{/�}/	g��~'�^vٞ��fjG��ãހ���9ⷾ��2ĵ|˫��ߘ����|�馛�C�7y��������Q����;�7_�p�	[Gt���M��sw:��y��7���G��g>�����}f�w��������Rj��7����_��9�u�u������f���k�e_@�K��F\�6�>l4p��R]�N�mO����O����8��Q���x�2���!�=� �8���y�M�-۞��W8$S��f5P��T���q绶3�7�� ,�Q@���c�r�Z�yZ�MЂ�F��[�:��I�G�t�x�LO�\��s� �(�����/Io�)�ލ�W��-~a:��h��4����_��Wm|b�~3�g��ވ(��!��]r:���L�ۑ3�1-��s�e�Q�7M��g��y�>�Y�;x^rP�g�#.q�W���u��0�Y�)>2t�i�k�Mi���*�8����jp&�����[��ҿ�?�s4[~|w)�����W�bd� ��#����.Ďu�
�G!�bCc"��2eo4�%�j����\��>��L,L5�W����o���9<^���d#g粞x���x�?f%�b�-�QМ<R� S�PT��NFE�*��p]�-�;:����L��>z��_��g_���}	GQI�.7Kv��	�щ6�ӸAH3|��}v#�ma�SU.	���6X��G����pl��+.t7�K?n5<��
���,�u=�댻��K��2$�
~�%���;k��2�}�]Z#�w�yk:�V#c��݌�Sʾ�{�7}�S�*E�����Ou,>����Ks���̀��!���E!��t��O<^����1S �@��җ�T���K"�%���������o��jF�_���{��gyֵ�]]���G�������.����Б�7^��P�h��,���@����<��35�픧7]_����{bz��ǫsc�ɋ/���É��g��o_)�cIٻ�/���:x��>�+����k���}w�1b-~O�7���q���]�\�i�_+o+ǣ�'ù��[�k�h쥜\@[�|�_ફ��t ���.��gn�e��!��?��ӻQ
���ʷ��A=�h4����'q�'��������[����?����'?q�����%���U�K�$�ǟxl:�Y��^x~������	e)m�S9��[���C=�c:ON�/�x������-��g>Sy'�����韦����~���|��$C�\}��$����82�
�:�=<�r��IG�e��t�-��~�%_�����(3:�f��O|h��,�3�u�	{c�Z��of��7wx�xo^�������w�����ۍ?�%>�J��|'� ���K�'s����g��x���n3���4�����\҆��V�a+��0�ϯN?f���m��G��Q�®�/}����7�p�U�cp�c�X��M7�L���s�G���w�K���h����i찾;�d��x���$ȓ�#m|��Χo����׾�����~��8�5�����5�*�9�
�����ۻ��?������s O[v�ߝo�)�K���gΧv+��Y�h��a��7�΍0�������"���Q������HƠ+"XQ6���~�>b��]8[(�D0�S|p6�؍{k�#�K��+Ȋ��|bmS�e	������뤨�YaN���lR8�H�B������K�J_��n�K�?�q��A�n�ru����q�J��u��c ��.͒��Y�V���ڤ{G)
�[������t&��̒�̩ጭ�)-�K��fi7�uZD��}��W����\E�u��k��a��ؿp��E����K_9��;���cW�/��"���U�Q����/�ѿ(J�K��9�B@�w�}��8�ه�#��OGq�(~��ߟ���L�d�����R�>����h.���k�ɩRW֞����oO: dݦ�?��?�������?,C�  @ IDAT�} ��+�Pv�ĥK/��:<�x��%ИZj����z�F�o���Ug���S5;��o~���i�����n<����1J� #@ܿ�(�W�2�Գ�L��~+���JNJ�0#�'ߙ���鎋�Vg�̄2j�����D��넢=9�F݂w�&��R�s��!�CfT�Gy�CQ�\��)�%�1`�{����W�}�f�(��疛n�`��)�v_4nאS\���D���c�+��������o�f��x��$���ϴ��Ǎ�y0�`�P>���K<fD�jSN1��޻��3=���%zq:�c��]�r��S��s��o�������Ͼ�wS�Z����[�A�6y�cn���(�wM����k&�B�m7�><5���A�ٍ���Њ��m:o|;]�:t
�c����8|}���_��8�']��t��Ӑ�_��f��z��Z$��;q�߷w~s��p��渖��|,�n�؝>v�����Mw��Y*x�/�*^StN-_a�{�%ܺ|���y���kڛ�����LV�8�eŧ��8w��L�M��}c�U�s$�K��B�����Ͻq���������<�����/=K����G�4(h�
��>F®�,h������m��nN*�g�T�!����̚#��{�f���%��[����E�qk�a��#���@���{��|���u'�gu=����d��<5@Eza�����R#��$>�#eҷp��m$���]�Z��%����\c�r�8�gaNE�酷�bk�L#�-��n@�I�:^M��k��Xw�@��hZ�覰�3��ƳA���1�0��r��Wp�^�;{��@���A��Co��ˆ�Jz?������	���QQ�{*C�t�������ij�I��֕x_�)X�9l츗�������xoZ6�g�̠$���g['�0���[;��ؙ}Qr�ey�;��M�B؁��K����馭ӭ�ܞ���s��t#`)G+����t���x��R�����������Lo�A{�t�7�-#�ָϬ�%'	�������͔�~���t���I�d��7�S�r|�N�_��_�������P���;n�΁�9�^=��N#��ޚ��p���X�D�vd��})?�����/D	��\� _�v=��Yg�}G�ȩ�#���������{�ߩ�S-�)}�(�RF���|�C������Dd��KN��:��6~J��Geǉ��x(�2����Mf���\�U�7���ϜL�ޑ���Q��0yRm�]������IVU&B�twY��E��?^���'KG��Z�~i���>?]vɞ���R'r�c�w�X~e F��A Ǣ�nN:��ɟ�2��j��ʑÇ��}b:m���U30��K3w�:�����Sǫ��e`ulB/ÿ��TK��1�i��b0j\�vu:ז	^�oo��Y^�(��N3�:x��ٲc�t�5WFo.�ʷ�[ؕ�3h�;�1��K��2,���J�����҇���2ڎ���+��f*��<��o[�o:��_8K!�P�{�.^9��܌��� g�����%}����4�#�K0��׈M�x6n�^����=h5(���|��F�N�oa�!�AR�ύ9���C>��)���m
8O��@���K����n᷎K�uO�����5��^��zҩ@ýhH�Y���eE(^a:m�tX��m�{>�id��E�":0�H��������ϯǁ�a@+ϓ_��+�.�7:����z}�O�<���Fl����ˣrx��*)�_&�����<���)���ޜB��d
^*�4��S"�;��yK�8�޹�6�m�z��Q�C�t�p�NwP���-pu�@�N�\\&�;¬]F�R��S��$�5�fΟ?�O�0z��|��i����%WҜ8OgI:O�)9��Ƚ��o\>��Q�JAc*�d�b�h���l��tⒸ�
���:���FXR8������p�m*۴��	�t,�BK�8�W�"VH��Ar	��dT�l�0ES�f��S�FgK4�훲�.�K�O��B��O���jf�2M\�0�C��7��)�j���-LK���U�3��9 ɮt3|�l�Q6�Z��O�$N_c�(�?Q<(���Jsd8�����i����춭��T~񋧲g��3��r�]�Yˇn��@��r��Y��*�Njrd���w����~>w3�_��޵T!d�L����<��N��Ͻp0��������D�}:a�ԭЏ=�x)���8
�U�٘�o��Z~c	�E�x�����0�;�QD��~e�x����^���k����ޞ����O�7e����i�2o*&������c���v�,^��.����/g�>1]�{O�q����[r�#>���H�cg���cU&�o�ۙ�蒣��m��Y�d�>�Vޝ[�+�:f�B��I��� ��ꎚ���=8�đ��6��9ߓ�dGt6�A�RWU��9Qzj�\�-���J��h��]N�w��s�Fvwʕx��Y#⨼Ů�m@Cl���٩]����F�ݴ|�4�Y�8)��sφ�i~����O����CJ�N��K/�G�^ti����e^��ґ̱�!_���Y7>�_�f�jN���0��7�w��������#+��2��%��hn�>��q4\�N��ि�2� �c�akey��b�uex`\}���R6�?��ӑ�q㸺P����:	ʒ{i����N٫�L]�z�XVx?��:�e}�˽�y8�z9��.Ίw���#��|��"��P";�jIz�mꔒ��{���5=�5�Yх
wȭ%`���0����0�����7���������T�վ#�Ҋǖ����&���y&�	��n%�\?��W������~p���z��Б>4�m����wC����q�;�yy����x\RI	�'e��z�h�>ORu��gqu^;�pA���>-K}�^�OG˞�S�i�&�=��u6��������Q2�<��t�DxO%s'D�'��y2�n�Vf�J�>u�奣}7��5�:ϥ��lk��4H3�lޔ�C��u[��A����)��3A� �6�s^5_��v6�.�Xnx�����Q��M�R���dR�Ǩ�9ޱd�&�*�&�_�h�ա����#���(/��j�Ӳ 
�x���������O%J�$�$�J)�E_
 ��tgG#16���ϲ2�ϟ� )'���4��=�:�Էp|͛%?ڍ?�6�}��i�a�{�Y{Yp��L�5���q^�a�g�b��Hvxvb��8_�u��8 -q˟ �4ů���׶�.0����m4K�%ݍ�����F?nұĵtkwv?�۔�)��Z�0�y��Z��!��j&�����]]�%>�Mwg������/�6�UC3�o�x,��_�B^���
��(CF.�H���
8i���u���%o��z�B�xj�I;���}���1
}.����ثQ\��2:�co�w�+ܡ5ɭw�* �G�+���{Wn�Ng��ni��w߫�#�������oeo�S�(2fK�a��qs8>��w)a�Q�x����7t�ֹ%��5�\`��~�d�#���U9xe��)������n����VN�z:=�`_����I�z�&��u1��ш��2�1���dxr(|5��#��i��c�ރ7�e�%u_���k���i#�M��ݙ���׿6},Ǹj`\P� ���ک{��t��������C�Xf��+3�)���R�/�1{q��)?R3w����kkR[�%}M��J�&y�tx�\�y�����Й(/�{fS���O9y(3&O>^�{�N_q�o#il��L�ݛ�7�w��I�襠>8;}3��y�9�?8�g��Qiλ��|�,z�Qn���������u�:=�5݂�Ep~V�f����,�����vk{Fu���g�m ~E[�6`�a���_�m~���}�G�]��L�0�{y�{�X^y:<�~�׳�!9Q�|ᖴt���)g�㧽4���GҲ4��ݪ=�8�xX����Nů���H��%~�hn����ͻ�;}q�Zy�:�������q���#�2��z��E�RH�B����}c,Z��2�/�:ù�\x~H�p[~���L!@x�}�M�%d���>8+-뺿Q�or�a�����*�yo�]� d?��.7��R�Nn�h����VqVZR9t)����(w��?~[z�TfL��N?������|۰�oOWb��pl�l��?Ҽ���-M�r��Ŀ����;L�aԍ���O�u�9��OAl������l�N�����I:�Չ2�=�Sq�;j�HNu�de�'x2
x�l�o��w�WJ#<�'��MgN��{s�����,�U
�����s��q,J�/9n�ՙ�ԧ>Y��o���(�gJ����.��ʾ���sY2r׬\S��q��ۍF���-o��AQ���9=n&�[Ip���)4��n�V�9�2#�r�fV����\�g�*`�J�ԩ�ſVrF�b��2:f�Z�JQ+��x�r'�?.��7�ɲ����g��*��+N�W�m�wmZn�)؄S~��_?������`z+w�X�d���eFw�q�t�=w���	��Ȋ�e5��M�h=����x.{^��RL�A��#��).y�x'N����¿}��/L�����s�����t�-���];]u�u���?\���!�+?҉�޼M�U�w��WN�LFdvck�β�Ȩ�wj��|p8���ATxtT�"�%y\3�I����#�ě@����������GՉ���/f����t��	o�]��h�κ�Uql<�n�1�~/܉�w�97�m{�S~����O牍>Oeha�� eǱ��o�-M��p)7:��t�H��n��V���`��qӃ�EG�*>uZA�n��n�	dڭ����7e��T��?B��S�`/M���g
�^�h���}Ļ�S�	K�=�p�<_��^�qu;ك�dۃMlaG�3�:_�|_�UQ�Ϡ�ef�z�e��D3ɻ��r��:깑_��5��ִ�?������9���#8�!3��n�xo���2�{*�9O�����)z��#��� ���7}_+�b[�l}C�,��:�զ���3\Ѝ߿�o�;'��,A	є�Z��)@ED�Of4L��.xCp�nb�Q���X&�T(	�P��Wqi~e������+�6��h�ߦ�gY�wS����	M�t��%�ƹ������5��Ì
H|M�{��a��0�4�*�R*�V��g�]�����x!����/���f_(L��A�K�Ky�f��v;�5�������0�A��Hë�n�愐u^YN���cg����چ���G��˿�;�}�f9й��+���=�M7�ze��_����%~J����Ѳ6^S`嗙�����������%�����|ݾ}[) [�M��y����;o׈�4y�F	u����ޞn�iP�mf�}ۣL*O�.����n�#��\�n�XQr�m"�C��W���@&��?iN'��T�+|�_4���Cn=�Ӷ�n�F_�*xa%����%f��_�*�*�N��[���3Ϧ#�Z�&�Ys {b�d	���8�/y����'�cv�n�ef5�)���R��uyܙ(�M=g��y��Z��<��Oy�4�q�K��t*�0n��E��=�No�Ț��m���b�м�(����;�{�Y�hg:ơI�I�W���&�V��=��;�G�E��eO��q������QKM*Bˎ䍴����-i���g1m�NgG����;�By���^��j��O4�|dc�w��^�V�8�Mô8�<i�2��+	 ���_t�t�����fI/���;Y�n��ܕc<��)�.�@���|��!�����Ha�uA����h[����N�K���Gz��S9ǳ��ô]q�Q��N�F��x�u������A���8G�����=x*M�1�1�k(K�>K�"eb��
3���v��e�p-�lƬic��:2u�e�d�lP���!0M?�W}w��y����|c�f���I�G���@�WX�rU���A/_�~��Ȼ!�CΈ{eǂ�1d5; n����{�B�~����]'%��{�5~Q�'D���YP{℥�?�5�hB{&�j�4c���
�����J�y�{��Q��
�G؍�F�C�`lWJm'�0i��!�BK4�)/I��j��d�3�u���q�t���&��{�po~.aڝ���yP�w�?��ec��n�
|U��^��
).�S0QH*�|���u��x���� �N����v!�����\�7^ܥC%l%���}2G�F���%58(h��0�̝nʶY��=�Y�j:۳��k�On�i�?3
Nձ,�H�5W_W��O��u��eW]��:~�3��:�s��}�E��H�9a�%t���@ȧ�Mʥ�K�^�/��ث��ۑ�o��V�[�e���t���
��J	eUY��������l�s���MO�a����ۂ�n��E�	���_��;<��)�c����3d�u�Nf]��dEwW��cW�x�+K�ݛM�w�y�tefF��{��7\u�YM���R�ʈ���wr�5�J��u��h�T~�q�d;/.\�eB-+�~x�5ft�=�eP�G]#ރ�qhE.��su*2��!�VY����%S�۲O�ʝ:5��-&��X���:':6q����qp���i�1{q{��4�ߌ�M�۶^���]r��M���맗�'H�����[Wu~8p�N��4K��_�B-�:~,3n9�@:��w��@d��Iו�7t��w��͋9����`��10F|K����.J� �&$c��?�l�v��t0��S�ߖ�i<`��t��k|��4�{��_�*E����<�p'h_��֜�3G�M�,���O��Ӗ��OG��puG��Np4;Nvǉ����֦�ma(�����(7q�q��]���x�a�����T�!
+����{�Xњ���0`��q�x��(��i��X3��6�s�]q&����'�����y�]X{?�������p�A#:�7�+΄%x�#�e�F�tP�$x��\k��/�6����aڽ�}7������p Ҝ�p�B�[Ъ���0�Iƙ��d�Ϋ�X�T�b�g(�[ �>��պ����N���G�K��Q�MQ���trgV�GW�-��vB&mH�*<�<����í�Ô�e��ҴXw�1�(�*��NgՆ���D3f���hL�]�w�گ+�]��郭����,qрU9���
W�1��\�aw��ۯC,����%����ķ|oxn�ki.��[�[��]rX�:0�3:Nuɝe�E�t�)K6�i��ht8{,�h_����ќ�[=�΄وG~��y೟����\[�x�Mu��ŗ����g�{�F��}�>��RR����£q��3 ���Y�u:��R�ҏv�hC���#���?�����(ZQ�-K�_b_�Aǘ�M�8y�q;�%::2��8P������Rh�����=O=�LuLЮ�AIU�ᗰ�l6����,~�aK�.�loݛ�Mg���,ug���׀r�Ã/NS�a�������.�W����r�j���y��d���eF������w԰K�������W���m�UJӚ��Q�":$p��L�N��8�3�"[�j�I'�K���Y*e ���	4v�4���?��|������Ŀ���Uu*� ~��y套G���j�7��_O?��#��-�?�͌��H��)U;�����Y0[�Hc����we:(�M�a�;3������ȝW��q�&���d����!������~�����>S��t0��M�o���1��j��V~��*����dUo�l�!C~��.��O��?�6�[�w؆e�בH�k�7�,Sa{ʤ^a�s�w�W��&҅/�Ř�P� ���F������ށ_��J ���恼X~��g���/��3x2�2���[��k�o������W����k��;|�qX�k8~�p��e�;,��6�>�`�|����h3�h<"��ͼ>9ޖ|~��t��b�"��]v���f�H��#6{G�rZM�Ƒg`�oS�sV�{�9g3�`�7|w�ḃi��n�p�n\��ۡ&�;�����Ɓ���u!�9��7�7.��80���4�Y9�o�b�a��
G��C3��Y85��U�W4i\RR����i(4�a+:0�:���PnU��X+��{�wر�c$|�/<��7"o��ް�G���0��'������0#���?ï�����M�M��g��V��ƥW~���-�����4Jg��Ka�Pq���io����;�v�\���]���;l��~!�p��Ƴ�m�%����M -�ٝ%u�*E���c� RloH��Fhav_�sڛ��p=���9%�u^z���E��(�
��ΜBf~E��G��ތ�:m��b�^s���/~i�+��Q$��������+7Je2(J\F��A��k�+����,���]Wg�k_��R2E7TSҏd��): ��[��賂PXF�7������6�($Q�n���s�}�h;�2@�<�L=�������ߔR��~%G��~��H�={.���_�U���M�q������}u��x)B���)U���F�S��z�m�唪�*���W���U�ɬ�cGs�Pf	�����5Oɳy���Oʻ�W��2������|N�K�ϩP�-����R���^'_Y�4fJO��`C��L֖y��F�),xC��y��M�ǘU�:F}�SZ��g9�M�7G����;�0��U��$�wh�:ǩ�{���ҩ�ū���U��=����^I\c_��yi�:ZG�̐�����$�d:}���ģ����7#��U'ϲ<�7,�<�q"��Xtg�W�?�(>�izQ�)W����J��^�_����p��$��,�Ny�n#�f�<�B%��o4�;�e~6,��f�����H�+\l�+�U�F���h;���[���n��~��PFħ�xt �^���ңSn����Jٓx�-a
w�UؐϦi����/�7�d��A�K.���w{���}x?@��&���|3x�����|�������i_[���6��_��U���h
��^��D��kn����ё�t�4V:�?<��c��9Z���Siʻ���Ð]~����Σ��W���k��ti5��E��̇�<-9	Zy!���:l�d��U����3|- �<��
X���~JP#��hc|EÜ �!��+7�� �Á�V=��?��Tυ�
Z
�ў��n�
m'��[�����ܤ�
bln�Y���Ǩ����O�-��Oǫ��0ܚN�����]��푆�M<j��"m⒞�ؽI��Y��7xq��ͯ��6>���]��]�2K?��,��hz��ޗ�#��c�F�,���K��F�.������+9���
l�����P���j���8=�K�~��ڠ�)�p�n)~9J�5�Aђ�Ͽ�bmp~��'�g�{�:tGϛ9��7���,:QK����J��{@y0�����N{��u:#Δ��+�y����t��}��\�r���;1=�M�i+ø���}h"���#ݖ%}�{߫�����ʝ7ߚNQ���w����`N��Yu��v(��؛q���*>����VPx~��(d�b?:�u�ݫ[�)���{S.�5�KS�ƚ^x��^�g�y�I0r�M~�Y�[9!�qLE2�Iv�ĭ��c��~p�(�UV�����Ԧ���RO�.�Iۛټ�r�UP�k�(�2K�\���;�UxG������c�<������zq\l49Ո<�������:�pm:�Q���M�N��d��Ν?��u6V�nα�υ��z;*�:5Y2�·*�����S�}"#���N�9��,С�T{ln���tX�?���G>9��Ȼc�4Z-Eۑ}���������<�Q42�[ܕ/3���	�?�([ݫ!m�'���#�ֲf����î�����5l���w!�[�s'�L��z�[�����G�s�O��<ӎ��
�o���C3~:��u8�ڔ?~�hJ|����~�3�^ȴ���|�N��^Î78�I�p;��c	�ćʦ	��w���Ӧ�yg/���gw�o��y�2]q7-fb*\�;�2�i��[��jb��i��f��u�
���y�7�����oj�w���.����eoN`<�{+؏~~w����W0^(/~���)ۨ��0*�h�hX5�ӻQ�l�JkW��ѱ��4^�.*�?Ϻ'�� c*0��9���m۲�3OVe��`R S��I|
̮];�=��v�x�~$tn��<������� n[��Ƽ�ǧ]9K9)��_*C�s�oH׌N\��i�l�ؾ#�rFa�zթ��L��r�38�<'���}�	�N=��ڨ��*d��p�4��Sȶ�����~�D�-W�]h(dUA�J^^ț�?p��2�Q�y�_P'=�����o�G9)|��6rSF5k�'�W�x�o��������/n6u�K�	��Js��M���\zao:�{�{�Sf4>d,z�
w��w�U!���� q�W�4�{=�0F\��հ�9�pδwk�KAC�1����>;�� ��e6��#Sŗ��Ol�tF�
__)+)?n�~��G�Wsk�%<�HG��
ҷ{SND�}��{9�����ߪ|�y������qh��z�F�5��:��H��|�q���̳/M/$�?^�ӚٝͯG�����<� T�?�T�8<S
�,9A���J���7����oK#��m$�9�ѡ��>��~QN���(�O?�B-�8p�@-�B�Mگe�ۻ��(�;�0>���x�9��6����[�W����W_~ez��w�����'������˹��IQ����D�B�����y$o������vG��K�*ד�L .����"i�w])� �2y�Wq��*�N��e/�Eߦ�����ـ��f#~f���#?{xz,��gN���3���3��9�HYGmӡ�rř��p#���%�
�F������g�����1���y9�<~��wx:��w����g^xq�/~+؄��m���zz��_NO��L�;n�|�I4§\�W��tK�NF��G���r�O`aq��<ඞJt�W?�_�5����?�{;²J��"h�
����g&�xC@��m��U��t���C�8�lu؀��$���a��3�U��O�A��=��l�z������V����S�~讽(�E�I����������R�,��)t��fwe����n��s�ɛ9��CI��цD6�^OɼX�<�Ã�[�Ч�4���:ox�=WaN����Y~�rP����,���44�5O�٩�g�`穼;�okNK�wX7F���(-������fV+c�5��\<Kީ�N~n��	uYH;mƶ�a{-��]�<��/���뜙̹=�N2ҮL�Dr�M�?:����A�N�ݞz*iu�P�-s}H'۴9eE�(��H�^���S7|CG���w�sk��ߔ!��ӡ���]`Y��#��B�G�w� >k�� ��{�X���.α�y/���e�O}�Z�����M�2���T8�KSe
��B���1��撗6���&U���
ʕ��z{'��P�� ���L.���U�j�sjȀB:*���s�ll�z�L���ML�V�b�#���TV��87?��B�$2'�d� �ح���홹���a��>7��Ί&���G�L�Nŭ!��n^� ���x}w�e��rӧQ_��M�j�Ux���D;�2�;��?����d����Ba�57+gT�N�ټsz9J�Qa#�:�r������Fm��#qR��)�i&a[/�����C1��4��+���}�K�ؕ����o���M���֥;�)�§���X�\m����L`yMƭgt:OD�Of�|ے��B�ҙ��{��v�-��ru���5���x������7�G#�|��|Iw�X�O1'7��*{̑�h�c�[�.n`^�"/N����;�F����
�#�잃g�9�mfAJ�%a=�Pd�����J��̖N�)N4(C�B�j?A�*O���7��j�J+#�m(ܾ��8|��phH�@4�:�op-o�]�a�eAz�/?y��w���ӏ��'�dʋ���H�+�G��Һ�؇���H���,ij��(�[�e_��������_h9�q����fi�%W9����^�l�t�%�-[7�(χ�W�?��q����l��g�0�G}�4?�#?�VC��U�? ;��5�Ƈ&1�{iڿ���n��;���mnL��sk�x�/�v���#mP��q��|��=���Kg�N���vz>���+�Q��eʷ��'�!~��ۃwܘ�}&���}3���-��p��q,�T�y���f7���e���pA|���~4tI�=�Ȇ.P���̇W'l�<�U�*md�;X�D~ר��8چ�Q/�K�\>�9�t:�n��ꃊ�sU�9�7�:�2.��i�|�������tw|�<F��}d~w�����>���ݶX��c�����Yu(�_��2��2؍�Q�l7���p�</?�r�ƞ����]+� � x�r36�Ɣ0u"N�v�S
A*�MQj�g�Rf4o����(��n�R�*݉��&v6=o6����*��?sƹ�q
~�O%�~�jIJ�9���chS�'��T�x[h8U#*�Q���F�gw��%Ng�&��P=(nQn���,�]�~�]�������ti\6�)�\�'�o~%$0�R����xz���!'=�B�6�bX'�D)�����b��U�qoC�P����ʊ_���� �iw�%%+�ƌ��qQH�|ڈ׷ޥ%H����Y��#��[�V0�栐^Q�W�	�-#N'��slq�V���Wv��#��|E���q*%����=�*��p2kЅmwf��k|��n�c���P��j<c��l��N&��SFX�cd�id����HҼzo\b'='3Z�2�[����͑�=+@��~p3ہi�ܟ!�f�ԩw+<Ń0�R��D>:;����6q��ӳ�E��'���0��8�� `*o�^�1qO+EZ��Wx�f'��	��o��wǷ��3�1�^ɬ�v_��N��! ��T�'���믿Y3�������<�Vq� ƺ|�o|�ik�|o
�v�
˖���ȏ�T�������gG�[�^d�\�VG��2�����|哬lϞe"�S��s�WGn
�C���2�-q\��N'��+�JP#�z|et*�;40���1�G��_�[&�L����ǜg�Gn�;���z�����}V�[zt���k�Rh�@�4#@���h"3� itb���.3�%�=��V��X�Un��v,|�&��G�m��ܚ�����n���/ߗ�+L�x�4��`�l�>�H[���iJVy��;<�Y4��]=�<v8i���EJ�������~���,��]� ��N��HE;�kB"xu4�4K�����q���C?��1�Nc9�nh�o�Mg]��vQ���"r�W%��?��8�����b�:f=�����B"�F��+e@䎜���fּྐ���J�S�2�cI�����V�g�w*B�U�Fr���KcP��QRg��!2�f����fSusa@ϖ4�����otZ|<K9������̖�;�H�9���M뮣=g�X����8"q6�ըq%_͕a
�P)/
�ǈ����L�0�
��#�U�c�����)�t�yę
+iO_�D�j*y�NG�*��Ǵ_x,�8�.��,A@Ö(��q������0:�s����.ˠ��5�/�T�����pp���(�{)W��;�歸�uzϑ��g喠�7�NGşF�7eN�AL�����HGi�U�/)�K��LܱcF�ӱ�|[/*��G )7�R�W��m����SH�w��%��4O8�D��dz��S�sqA��p��Dl�;�$���)W����O2��a:k[t��4���*�t�Gˬ��^���F��
�#a=]&(7�p��F���B��4�;�H�f�x�N��4����ҷ��+M2)�ˡwx|�ɴ]�P�]����i�:	?�X�7>y������ܒroV��充gȗp�nR���i���4@~:|���}'��X&����Tb��ɔo��F�9�C8n�#�J�&����O��f6�p�3����S�� 3�#꬏򅆸V	��X�Xќ0�B+:��[�+�L�w��+��B+�;%���A�����Fg���)^ő`�7=�w�r�u�^����1K��pO�g�����N�w*��+�2��7���dt|��];2���{#�Y	yo��l�䇲�n�z�e��������������v[�]�o��A�MG�k��p-�������ٴƵ�n�g`4��n�K�<Z�z:�x{�;b��
>���wt�K�\�+����3X:\��(�5#�7K�jiq�_����}��F�1@�ne؃���H�m4���<�̷M�c��j�t*�[\x�~)�����h�]����('�{��e�q�	�vW�oxC�Rf$����c��=�Wf$R H�о�k��|��.5HJ���J�����a2"22��Ẋ�V�Y�	��H<72_����ϦQ�j�
f�1q�����o� �_�e�ʶ���
�sr�	ޓ	�tm� �_�v+�3lx�����ٿ���QB�]�^2����)�{hV_�E�������^�Q���k�w��}�cN���F�a&3Y�yz=O*�];}�G�I�̋���J?��yg0w�F �ܱ� #o�T��94�S� �w<8xn�n�:��E/��1��.��ɒ�Z�Gk�r�#��r&t��Kx�{�I��J���6���+��c�����'�R�w���1&�� U�|0��$p]w����~��2�:���5roz��_7�UfOǙ���v5�r#\ʮ�e�{xK߹�'q�j���G>���T�v2�ǔ�N���Qt��keG����i��8~X´�90r���w��MZ~�vi�k�C^��_�~���_ipkga������;8}�@D礞m���3�=�~�K��D���n�ʜ�rS�u+�d�j�Re��%��oOh�%�
��Uz�Шnc������;Ĥlt~`V��Uov��#p��!6Џ�.i��
KK'��y�r��gn�Is����K�%��~=2��|�̕�$k'K�e#�ߧ �o�p��WF��h�H�q��''k��֎��&}�`����w�	T�j���9s�c���,�2��4�֤�6��58kK�N��W&9���m�$�4�| ni�͢��t2w?�+Ξv�\����R���*{`W7����`�)*�;x\��N8�Pڗle�l��p��c���<�ک)_uQ�uU^&��7�mQ�L�r��S�I�,�-{V����y7s�kx�x��E8Wݲ�1ĩO�\��{�{��K�lv��~��{ӤG�MΕ^1���~��h��ˁ��?E����y����$��\K��%���V��s�%�j�I��ʳ`��Q��j<u�w���ПK�
W~����~��!ak�w����M���OZ����7�V�l����j�������|A��o%SYT����.����.��5S�Ӭ
�~z&>2�U �z�K��J(�k�B�pf����e�|�ƃ���2�����oz�p�U�2.��M�xo�g�����u�V�>�U9�=+�O���g��tx��񷇻���֑�l�Ȥ�a^R���äe�Dn�V�����[�E�2�����En�^L$�ˬ�͓B
�c�����wP8/5�.Q�}�ց�r��[G�F�c9���F
�h�i��戎<�)7<x&7ZV����u��� =p��ɏ�Z��%���l�ܠ�XGtn�y���an�f�]����.{����
"���^�&�㱯;k���x/��iv��'|�����蜲�[�	jJg�+n�t��p�>Oݸ��Mip�~�Ro�[*���ֈ�kۛ������E���U�n:K�mVY�.�W���yτ�K��I�l�ɤo��][�V�C�W�u�30�o��ނn�;�zor�V�ɶ	�O)���LV�����`�(��W9/�/=YgpM����Vm1�Ec�Z^����f����mO0�m  @ IDAT�{F>�ne�x��_���S�w%����7<}Z�y*�	!�u��{���܎[��O�{����4���%{cK���n��^�fG��DO/H��z�fn�  @߿Zlӭd�l}#������������<�E������~w��&�f����|�A��8�֦����Ӄ���pf\	�_��6�8�ȼ���a��C�\�'u���˧:p~Ĺֵ�T��o�s`���V]\������*�.\��z�~K?�����Yuա1���FLf�Є�r(3NzZ��'��Fz��#�]{��ǹ�׵v��+?������\��n�K�j���Z��ֶ-wmE�FCނs]c�4��@%�q��:�8�#{�z�b���ԥ�-w����r*��%�Y��&�4���Y_ޥ����/~�˜��3���,��{ۀm�|��P�ЗW�=�����sd���_����p*��������-�2)�x[7�eݼ��h�D~�:Cp������������S9V�Y���O)>��a�_��s�\+��S�tLNo���)�U|�2o��g��6���L����8h��/�h՝��}�R���~��燳����_�f�97ߗ^mi��'9��K����ٜe��E򍛁�/�ۯs�����u�l���΍m��:�hql�1�$�j�5$��-�����驌�I'�~_���2�9���c3nI�*������G�C/�Nkh���~�(��N'`�!����2����$-�OI�̖ltv��d�M�.>�v����=0�ɱ���3]���Np�b0�y�����$�4��z�^,��4g�'w:7|�/�#��6䃭]���t���p��(����GZz�8�T�趕7����xp`���L�R���1y�����^�x�T�o�oYx�r,�����'A��=:�
�̦)+t�c����ϟ�����x4ν7+���+2FN6���/�<_f��"~3{�_d�x-:[Y7��3/K�ib�?��zJZy7}�SN�>���R�n@<���M�i�Z �N\xd��4:ӻ�Mω��;��/��5A|Ɔxl���>9L�-&�k5w�z��gT�xGߡ�x���g�l��K��;t���4��mN>����w`R��܋L�}a�C�v�K���Y�#!��Tc�����L`c�h74|:I<v	����[�b)����m�I�ܲ]�.ma,�z�%
��za$/��%�[����c�P鏬�<�!�WWI�Y�F�C�Cs������|�����M�c�n�HȖk©�z�,/L��b�m��z��?g�S�_)���އ���+����f�ě��^���r�6�v&]�+�Ʀ)t�?����:6ч&=:��]W]�YxK��H<��S��;r�=�=�Bµl'vz�o�ǹ5m���U����u��U|MMV֘����%׵<�.�^|1�_���9Y�(��Gѯ\��W�8/�o�{�*gi����E�1[����{tG����)���v$�鿋�+
�a�j���՗�r���T�<ʶ��U8�j��`�-S��T�Ni�<ܿ�f>����K�*�G^��,=�Ǔ�� D#�'���|xK���}v�o�@����oϾr:Ef�9�N彟c)�c�"�H���A�f���t4��"K�$<����{��[��4�(�z�݉�u�Ȥ+mn��jg�&vv}��18�ح��ҽu��I3���K7��;���.]�����)��o�~�	�z��~^���yn�`�#e���8ʧ�x�52��ș� #C��)d��_7s�/�r�}��(�<�e7�)4W�ۉ	W�p|��W����..ۭ��խ�N|��Dˊ��ݼX�S��<��4�[�ieX �]t�l���=6�%���F�XD��{D�'�۶��A
9�޸���T�~�|gk�h`t�n�p�f������'�x����c�ɜ''V�mIs򝔁���Zn�Y���,7r�����3�T_9�����m=b����N٤�W��,���ih�]��w�� ����i:��틋%Y.ҾF����M��T�Sy�e3�LSi��'���&\�^�C��'��C�TCuR�l�K��8��'[�\=���(��v��E��λO�K�(�7)61�>S/c/������)�˭l�]�n�Ɋ��Б!qi���h��P�E�qJ����Ta�꧁�X8�a��G:٠<��EG��g&~MCGU�ބ�H�ݒ64ąV5����(w*�$�5����n:���=r8��.���8W:��Țr����G���}b�&>����׼�%�<
���>�gP�TW]^��_p豳�rㄛ窿1���*8�%}�-s
H;cG�����o�﹣�7>�:XN;��_�X�>�xx�������'�h����)��CeoZq���1��4Ďp[��K�]���+?耭k��u2*�<�7Y�ʣ���o�^��耗�:7mK���^��*���|k��}��\��%˩lȻ�oR֟���=2�a�?��đ�^��(��[�Zu��U�W���p��"ga]�?_�W����-���ԇ�vok������V�*���C�,y���إ��`r�49$�kݟE���{��>b�i+C#����o�N-�������vg0��t��қ�Kl?�W9S���}�w"� ��[o�9�������=�>{���7�<����9�8<��2w�����3��n�Q�e&m���&��.�y��w?�ܿ5���Ym3�0�b�9&s�	j,i��N��ίnG��l��og�G-�C6�[�.�y�F��Os���p�ɡ���=��
����|[=K�YG/�ȷRܽ��c[��Y��_^>����מ;X,?�"a���#��iP��K�ˣ�N=�	}0�mM NDy���o�~�ǔ�laR!�O�nf�����L����K����5}���-���^�<X~t���B&?2_<_Ǻ�E�z���2!/^ۂgՊ�o%��l���wiC���U9]ůM�X��Ev�����٧D"}��;wז+:�͓et�5`�`[O�A��o�<ܽ���B�wV�'���\7�ȷV��7�>�<MNy�%|��<F��:t��*�0z�n�|3��ݵ��'"������+���VGg'��+Y�{������$�=0�h���hM]K�I��K6p<��i��2��V��E-i���l�2�{�}6��1�̄�����cٞ��ʝ5�����)%<Mjne���ߞd���J��.N�LH�O���$�e��	��Q�z��c�%��W��L�Ok'��F����m�Nh�F�3A6=�9Ӓt�C�p�^�a�b�a�HC�Im�|K�,��'�F�uV�!�|#�\���Ed�xt����
�܏��3���{�Ih6������t�[�h|����!k�.p�L�;�?�՛~��-v�KZ7��i�Az�j��ϓ��6e˛>K���d�ץ��&��~S'G���ul�/�G�XYp�d4�d�Qg�c����"�K�gK^e���]q<�J�~}[g1(��k�u������S(�R.g���#=!|��$L�.�>�q�u����7S�G��	_8z<�#'ƍ�)O��W)ֽ�}��eq��H��DeAx�e�)[�i�q���,���c$���E7l���s}j'�R�&�s렒䇗LR�,ԭ#��?R���]���-m���]��_�y{+�P��x鳛!�a�+���>�˴�SA^�f4R&�������R\�����4��u\�Ql��Bu:��i�Q��tN[�jpn�^�v��L:�|#��$u_=����|a��_�A<̀M�~�s W]�o�a1K�3�r�zVN�X�|2ׄ�L��Y�τ<9�;'>��؏�u`���G��&�,h�w3�B�_:��t�h�]i���Y��͆�����wUz:�x��N��}ȴ�W_[��stܬk��?|�ËlC��)��y�r�`��4yt��H��6%a4ۉK��~�X��L˧���·�J�G�r���+|5?�<ۄBx&T:����<Y�����$��p<�V�gsp�'����WW�0ܦ�o�+\4��/ﯲuS��c{l�sO�B���'\Y�W�٭��άM����Ë����N�{�G:�|˽��ٗm�H���5o�(|�;�{:x�o�x��k��4�ӱ�u���і>�C󫗼:�p`x<��M~�S}�D���)x�T���I�P�h=����񥃾Ӄ�+x�Z`��#{�������Ǵ�ѧ�;�<II��������[��A�qDK7=u�����Y2�K���v��"/|���l4�K�%�0����d�䣏W����10�M�E�U��z�>\�9���9/P��/�ji73A-8���>Wy�Y���_�B���f1�k9�A�y��!������ȑ�����$�y)4}���r&)�DL�̶�LL���3���9H=y�m�N�,��ax>�����C�=��ß����V���O�E��'�F�W�-��M��u�"ǚ�΄Ȅ��[o^��n��Դ,�3V_g`�]����$�$���O>��r���^�ʈ�m�$��u$b������y2��~��g�ʫ��4��+��?�jھN�o�k�m�'J���W�kd�4D�N+WN��'�}?�W����y�%�l2TanɣǷJ�m:I��tR�8[n����|����o'�Z>����2ﯲ��,�E�tb�3��ց�u|f�>*�Ǜ�{f�t=��u0ܓLH��%oqtn;����
f�h'!?- 2�Y 9���#n�����Yt��Q���&^������|��\�8��Ѳ�ol��@�:~_�%�|q����k�o���l{�uґr�>�Ǧ���/�.��n�熳�Fe�}�����仡I�N�9@\�I����|��,ytX���O��axd�*�t�>��UxWi:<X8�rV�ڳ�IH��:� L�˱͑צ�Ȕ��u��bV���q#����eM�_����&�wn��:(�obDvDs�jA�P�:v+8x��X���RK?n���8e32��{�J\���y��;�\˥W��^�08t[�偫�/�6�V�G��뀑L���u�8���ʎ��éޮ{�-�<'M�n/q�O9��|y^�x�ҔFNN[!#g��k���rj���sʝG�<���[�+�|oa^�7!5~��\�O(lۡ�du�\i���,:��8�M+�\�2v ,����"Bm3�������Ko��VF��K�md�[\:=�	mi~�X���͎%���y�ϡ��-<48{�qdn���ɾ�Aڼ��Р����Go:��S4����ܶ�޼}~x3Uw���l��Zn|h��Fnꫮd���/�dG���}`�q��]m+�7�জ���x�+�g��|����"��j�{S��8pՅ���z����z�K�0������ٍpc��IF�k��V����m���!v\�Ӿr�	�,�]s(M��5DJ]�t:��%1��k���}@��Ld�m�g�1��u2ecK���]{��i��-� �Th���k��z���z]������3:�J9�gqߧ�IN>���h�}~����p�꺺۶���%8��"�A�� � �2�/.�V�ݣj��ki\V��=R�g֣P�s�1|��{�?�`�H}����/s�ٗ9��qN�y��[�ttʍ��&�/^����4|�gۉ��u�Z�a��������Gج�"׾����s�ۋ�p��)��uR��5�S�I�&O���u��+���y���1@�yV�����q-��������T2��[� Y�g/2�/��֗�u���M9z�k#�_�\��7.�;=��׎x�h\x��C?i|W����pڅ�/7<�*S�YE�3��'`�ҟ/77����-�Nol�衇/�hU�� �+/����H�Ө\�,<�C[:�ZŻa}XM�����m0����eV������B�i+7�>��HV�jKs�I��G��aSMp�WX>�����|<��W[����^����u��ߵ����]���ዻ��Ҩ,t)y����J������8{5\}��^�s����ƥ��oX���j���7����,�)�����n�̄����_�!o�;�e�E�&�q��|�E�C�VM��i�4��K�6H�El^���`1 �k��o��r{{�@/n��hH��\2����x�`��}�/��Lp�����rim�df���:d��E�FV�Kׄ��-c'�N�dؾj .�i���G,�M׽~`}���O�X>^��c�=y�>���s?Jy���9�9��y�!,���#ox$c�Z����mO��JIG��e����.�fd&ϵ}�W;K��	��������ٵ��wo�a3����Y2���g9H�V�}�7��ΝU%2��N}{����T�d��F�м�]�$�����L�r5q��䙞3�5	ǺG?�xz���FW���U�C�d��e�^i���ο��K����}��S��x��Q�^�yW�F~a�/��}�U��ŏߡ@Pi�Q��L^��o�v�3�	D�8{]=�v��w����?���y1�z:�'�
�mN-�����pVb�lf�N���_�H��I��;��Iz�{:���w&�Ԡ���y�x2'%]զ��\��\h�ܣ	WgzH�����`�O��G.�:4ЕǗ&�����!���x��#=��/=�^�ǯ��o��+MG-tֵ+5�`�P�9f@�����M�8+���U�������V$�Z57����dY��M)�(��:x>{�lu~sɆ&���I�'�q�19�6���4=T�n��t�*�)�./�+��F��W����_Ł�xhOk�վ�J���.�k ���ڢ��a˖5�\e����y��'+~#ߔ�iB�'*��W]m&���J��m��rj�<!�x�9t+[e//����[-�
�<����ѭ���҇�/�W�n�����º�����q-\i��}dm����|�3�����2��
���<g7ڶ��o�z�����������o���$��!�~z4=Y��<�v�����&SO"�ߪ��\�F.�lr�T��M�2��.�^�� ������m<�o�m�Onrt2 �ǯx�G7���(u����������G�$K�vr�u���Ǟt,��'%|�*�Xm�&�E��G�[9pc��ՙ�j�s?[�В׉ |�s�a��c@jB!M.��e�ؐC�G��o:�{�HWVZra]���	8�����v�|����	�/��������|�mz���oܛ+�%ӵ,V�����\�\�ܒ7̼���rx��7sO��1�7�{��~���:�]��y��Ý�?̣��I�eBp�Nޫ��"��1rm��r���޳�R��uɴ�ʏ�sh�&+�~��y�1`���4�84�����_��J����X1�_�wWd�������t�l�|זq���j���_���|_xMM�\:В�:e�z�@Wa~[|^��Q����UX�>�l���A��:�4N���x����ܔ����>����"M��ָ�?�yuDiW�k��aiD&-�z1ߞ���V�/�G����j������pVyu������w�ˣ�7��.���Z_��i�co=����b'��Ky�ǭ]�:az��P���*,��XX'�-^���\�.����]�e]i��C��L~a/^<2�׆ҧ�7}ě�7�97q�+~�Ay{{śV��%O�qˋ]ܨ�����
�qa��t�\#��ss�����h�0/���7Y�gs=�K]u̧��(�oT>���0etapd�K䒥?�X{�E���G�.x�-s����}������p]70#S`J�S����`�+�����a���5�U�W�<XNz�Ko����ɵ��U:>�u�K+���t�z���K�AK��	8���L O��'=���'|�k�����c���i�����_�G�S�.�����k����ȶ�ٍlq�s��[���C����F�KOނG�WW;�idIT:����g�BF������Z#�{�4<�G_/'�O�e��E�¬�b�y�_��/�dK/���ز=.���o��A��4[�8��pmy�M���ŀ�?X'�)��5ap�U�>kx���>G��=�,\X�ػʩ]ҿ}�rYO���ֿl�A<�����8��BI�J���?�'vqU�A_6�N�<qAO<����-���^���b{g((���N��;uw�Jp?p0��|�����s�<���6��}�?{�l�ˤ����p��'y_4��J�=�v���ny+'E޼�mdy��u�F�O��ڵ�2�smU٬6F�u��ӽV:����-���6��u�K����[������O=ʂDˆ�WY�+��U��u�:�}5�����]���UA 
#�Y�+��k��k3��T�R�=D9�J3]�x�6����fmG߹�p����X�d�,l�g'�Ph�k%1%��i����}���	��4�'9Qjd8��1���S8l�>�;|��Ra]O���z���^�*|<2Ks�Wp4vt��a��׫0��lG>��&#.���*�n,h/:����p�4�z�Ķ@e.,zK�e?7/g��䝼ڠ�8�h>�����iV8�R.p�D��-^��;�88��`�pꁰ�+�4�)���_���`/}��v��]uoɢу�l�{���Ţim�j��(�+�(������]^@${}a*�Y&��)GN�䆧-Q)���FVD/Bh�/T�x��x��Vn4�U�̠�y�Y���sn�V7����I��I�֕fe�ׅ��+ڵ!|�|q+��:#OZ��<��v��.]y{^`�'�qpu�t�p���5Mz�J�L�o�����fo�1����	 �ƀ��F]�W��h��a�]mұ�k@.o�p��9[�<y�ڿ�­�k/3x���r�pl�.�y�K}�\d��-�<����n��L��i�S:�!�ވ��5)�B���� s�K�.m���I��©��d`�rr�[��Pu3Gz;v�׮ӥ���;m>��	�����a������w�i����=�3�jK�s��Myf��ZN�k=�g�걒~��K���.���������5�Z[J~z�+��ǖ��B��y��z�����θ�俵�l&�q���gy�0[w�����~*��	��6x�����S'[O�_bQw�}ʨ���T,9~ӭ4L����$�c�y+�u����C��������vt~��ͱ������<%����ý<�Io�E�ؐmo���t�?��9
�I��9��vN����;��>x����N�rj��y��n����?8\�TK��6�6��	DmmS�(��/I���2��Tc���������9��>W]�/�?B�^�}�n��}�)����[m��6=&�r^e%|]i�6]��ʽ޷�N�����8�@L��p:����U�Wc�����;�B�ބ�H����sLZ����F:��Mc�پ���;�ڭPi���i7���ю1�<�H�豢�����V\G��t�4��) �A�؜aG���NZ�$�ma]W#�������TNO&������ঽ�[���z2+�VpҚ/�rDO����4����h������(l��*�4�]=�ܐ��b=�X_����Yr��T�uÛ;E������S�u�z�\¼=���,��~OssG�z4���sե<�·���{䕆0W���iF�tt��F�3�!^e�}�Ca�i�|xQo�@*���P}��j������
W>�;�Ն�֕�3(����W��PڗI�j��۪���6��	�x��s���Rw�.�2�C^eL��l��!��C�tě~5���!ˢ�p�?Z�
/�������∳ca�#�o~eo��Q[�vm�!��	-N��zm:��<���<J��h�������<����W]���� �)��/�����KG�N����䈵�vWʃ�8�U�r��΁���{aGeW8#�֞���:!OǕ1}��h̀=u�V���Oigad��l���#O��)��	r�4��e�y���y��������i�^�#�[]�n2�{��C�/3��$�	E�W�>.W����l�C�>�.ه�������`�$L�}_eU;�I{䞬��������ㄧ,�C�+7p���x�[ނV��WE��M+��5�=Z]���C�p���) '���a^v�}-H]d�F���e7)O�M���.���޻�B��[Hy0h�f����?|�����'�	e�v����S��>����?���_��'�7�~��a>��n>�{��s��R�oe&�*�u�޶E���'8�`K'�W�Կ�oe�����.��R��C�~ӵW�ΘMX6������4���U��I[-�ħueՇ+�*�w|)�d������oT0������V}3 �u��g0j������0z�He]:�Cx����f��\/�����{��k7�4��s-y�LˊtN{q����͖������t
o��r��Z���f:��[�g,}�ȹ�V��I�l{Bq=|��X��VNe�N�enYm�Hg3{pc'V8�P'�>:�,�sj����ԉs�d%�ߛ���-[A^�vˍ���@��I�a��'4��E�tx	���g�*q��ޑ+D w�Xɺ����W{�����~��D���)��Q����{dJ�!�0�#�<�]�r����[nnlY�����<���S�ƖY1\2�F���r���A��/�d�&.|�r��s3ܘ-o�q1�A��k2{�#gSOe���&V�j_�Xv^u�b�X���4�����k��E��[K�i	��l	�"_k�_��0X|������PG���H;|�,mg�	n�����kߕ� �K�uӖ'n�x+m�j֓G(>_[
J���R�*7YM�n�X�D�Vt4�g&����>f���=!���ՠ��MU9��t\��B]ƛ�v��Ό*�:���ʎ6��],��H~��������g�W�9�Y��#�����=z&_�*�yҳ�y�!�j����68�
=���������&�#kډդ�ˆ�c�U�6>})�6���B��~�x���v��y��ݴy�������llu|xOO�-e�A���ʹ//����~���<H*G-�`���r0@�B��Z��}	�QO�?�škI|���6�rtc����2L?S'-u=:�7�5i[�>�l��%�梫�i]�k�zj�4OY�pdFCދ�{���E�&����t���W�
�z�+}��i�>rV�C8W��H�2O���a�?ɶ��yWa�3���]�п��{���g�a�[t��-�4�V�����e�k��N;5a���{_M�����;5��N�p�s� )=����<�߱g���&�~�Ÿ��~���Srs/L;賋l�ʎ�o�7v�Ch�S��V�)����h{���Ϸ:�2Jb�1vL��x�hV��E��d�u�S/��Sx�_Z�ѓ|��Q����hW�d��2���/��Uat�z)�G��W��z�ү烗��:���w������^uM=3��}���?��p#�~�ɟ���,�~��|����������o��ȁ�{���ۓ$��l Zo�=���#�\�2��Ǥ�M}lp ~ϟ������6m�����C�z
;̽Ըu���۴�����ˤ����o�;b����*éK�P�����׿��|��i��=�G����C4m�����U?T-4^�ܟ\���ڟ(;u�36{�[��]�3��B����q��0]��ϳ�f��<7�X�b^�KG�QZX��ՠ�aiķl��ꐁu��u�t�K�s/[��|�^>��f&�p�j��L6��)2{����u��kL�!�<}Ꞧ4���n�������<�<��|<�����y��6\XXu���)���;�K>��M ?�,_װ�Ti���9�J�n����Z}���{�^��xq�`�2t����;�t����S�h�I^�0� [^���⊦0�����Vp�Wr	׋��-��h�r�.�u:�$�<^�_��=�h֕�xy���#.�>\����p�JC=&G�4^�Ӱ
�Wi)7>�r�/�O<L�� ��؆kG&�\{\��_x��D�v�����J/x�pe���P��ߟ_���q«&��P;�5PuK��? kîcNu��/gOC�@B��1�z.�׍��X{�N�����~����]�NuK��HX�fЩ�_[
��/m����Ծ��G����{��-.��,��c��.�9�.�ݪ���=�p��jK��@�/��[�#_|�
�4����ni�ӓq���Y6��r'������{to[a��~���U��+�r��NvA��9iS�R�#�f����^�O�������[�N=ɕ<u뽋�J�[_�ѥs�˧:7�	����ٟlr����[���J�z*O10�וk��������î�D=N���_�IN&�/3��u�f�{Y��]�r��G|��T��	>h��Yz�sW�*������l���<�u�<�~��8���>̫4?:|����?��.�����૯������ۿ?��>=���_��.�䶼��o�[���$��ngO�� m?-{�u�*�����X�u��1���d�"�<1�h���O���͙�S�n^����Yd���I=�{���yc&?DzVw<�x�27��qh�M3�>�"\��?���^^f{R�9=;Oc�Ħ3j��Q�º!Y!\2gk\����j�����I�a[8#����Yu����P�A'XC_܌�p���5�����\;o�F�6���ݤ�����t ٴ�yQX�'C��&٠���Fy��[��U�Wd�c�����U����3L�p`����S��KPk���ֱ��r9��.�Vu��Պ_�2Teҙw�V��1��șG��8��n�3����!�ő�� o���j*�ΞO�Nz`|9�E�a�7=�]m�-spV`]��+}7�q~l�`��U�x�}9i<��,,4^^`x�& ��7c��0�e/e�	Ei���yrȡ�upћ�������G��	��>yrа�zՖ������K]���
l�׶�kp�{����<�Y��h��{����s��U�K=[�=�l�����?�7|0�G�o���N�=��.�=�C���Z�Ss��0��2+��[�v�o9�rhYp�\�0-��>�"Y^��\���#���� ���j�]��G�N=X���1�Q� �?Oh�e�E����<�KN�M�uQ���˻�C��Vy�W����s�Y������He�D��ʔ����ci��N��j?�B������v�%+�e�������c��oF/��V��y�5��n���I9��F��^���n���� ��A�;Or�ף�:'�m'œ&O�	n�x��_N��Z#�����ȑc_v�pp�}�����m/t<�w���b�փ����/??��˯�d%�����c�-���	����R�/[����-̺�,����-��-�WDg<�^�.�Ν��>�����ß���>��Ù�v���T�ZG��f�����������??�◟��g!`�����-��Ƿm�u����ܿ Ĺ�y�w�n���2���bb���,;ĩ�K�q����߈b�{��QN#rTA4D�?���K���+��_���|��-���� 2�f��$7*��[�T~ݔ@F~^Z5S�֥d_�dwʂ-0&��0����ʡ�J�����O�zv�3�Kz�9��Nnu��C�U૳�#]GVXW�'���嵲����*�se��OG{�k�+�:��G��Q>��$��v3v��|�xr��r��>����GYC/�<�qh���_�X��m����h�O���;'��Ȟd,�'z�,�<?�`�PԦp���i�	fxG&q0�W��`�ӡ�� W�[|Np��._w��W�:�N��
��)�kӪ[��*�K�[7��BO���)O��sMzi�m"mɳ&��l_~�8[U�nj�li�I�\�6k:�p����-�ғǹN��|}��-O?�ޜt���eR?�/y�X�Z/�U��7�t����+�wh�
�ax���)�����K``'�Pe�Ǘlk"��y2����$G��X�����ga �e����V�{�-�� �|��RҲ'M�r�<ۿ�����y\��rh5�|��KW��g��}Ny���^<�O�frp���j��F����=���UN�
�{�FSz�l*�U'ޢ9��`~y�=�.&����ԣ�,W[��<�<\/�͢"<��F�q�����e���|<��	��һ��I�ߊ�g,�h�(n�-oy�Z����p��j�K:%m&��%�H'P�>��aN���g�:��o���~���Y}�֫�E�̬~j�?�^�#��4��������w�����U:�k�1w���Ï���_��_��_������;[��Ex}�q�͎��3����m�;w>8��A>���;�7ߺ�1��?��_��>J��^/Hys�.YV�m}_�,���U��'" ��9/BϾ�L��G2����߿���?:��||�$/}�ᇇ;�@�J8�G�7��8��Q�`��ç�����_|v�������"�8�iAf:����T7J�U�5��Qz�!K��Γ�و��ɜ�p7��,e�Y`F�W�юm:�1-C�)��e��A­��0�Ԗ��CV/�I��τ7�#�&]!R�诎�Ew�\���&o�)n;� y��I�r�LpȁN�Ɓ�{�*_���s�oɹ�抣�����|i>,v��$C�#���0Y��3v� n}�|}Lm�BN� '<+D[g�C�}�������+fo�ƥ��G��H����tJl��o�\e�^|��{��Z�ܘ?��)�t���hܢ����T:8��o}/�М��mO�&^d�����u��ߟI��+�����r�Z��3��O0���F�}[N�F�����>�<�iuAC:�3�����+<�eid�ތ-��+�>��+C,?�F�uu�SY���ܺ�$��nxk;���O�M���J=��y��x2,ޫ�T�9�"�]	o��_�\�w��ot�=@xq��s����_Z�n'����-��*md�uOOZ�5�����N¥���|�g�ܳ��.�H��G��)�x�w��GmWN�qidg�D�n�8�c�{���dN����{�mP��4k�h>���d"���up9[�p+�߻��]2���ٰ4��b'�����Ɨ�0�ϩ��q	zh������9z�.��z�W���Zp<��N`~��U��1�g����û�y������`��V�㼗J#��|��W�_~���yJ��;o�G�:����-���Z^hWt���f��ˣW��s�V�7}t����_~����X��l}ZO�ڦ��z�s&�7r�·�>Ȼwo�^J߽��w�(�m�_����ނ�w�:�F۽'-Gp�V���Z�_[�"g��T�tx�L�Z��o>��{����'y��9}2ǔQ�Y^t2k��`K�iŗ��f_��y����?�������o>�r�6��<��*��A��:�tF�tƚk�=̇�y4��o����0t����x�59��Y����o~�OۑȎ&ϵ�����n>M����+ ;�w퍦7;���9��J���km >C�#y�z*���ޕ��M����N���K�4�Y�#Wʨ�_:��`�kpS���6X.;����VR����I�w>j8�i��7�	|xo6��W^��5�<��\t�%�p���~��Wxt��j4ʿr5����֭� �p<'ݢW�L<��F�������N<8�`�C��g �A����E~%[���+0��ax��M��^��e�%K�*� �2�/����*'�p�қ�8�I��{z$��8�r���9t��]ZÕgl��aQ=��	�;�~��������r(T�.T�ҕ9�:�EPNun/c'�x�S�w�Cۆ��Qѿ���Y�`/�=i�NzOQ��<��ƽ*ò�d���֎M�ǣ�w��+�0׫pyhḻ��UΫ�s�z�À�7x�4�o�<�&�p]���pŗ�-o��;Z�p��'�)�to���E&sHB
�ޗ^�]�&�A9y�{�diE�;��  @ IDAT��Y���i�夳�'�!8^}��s)@�,|�C�}��)?�AC�+.�y �=>q\�74�Sy�M:?��V�.�>��~f���N�%0�xi7�a^����og�5�&�Pl��A��B294�W@�׆3K+W�,�IeI���1Z9�Lqc�soTIJej�8R1se�p�ޘ{�"n�����n�չ9��>7�ǯ�����+v�P�/s���gՖ�!��wB
a�vBh-<�.D�z����h7���p�HlT�Gk�L����J���9��5���(�G����q� Ӽ��$��j3r�ɟ�R18�[-��Md��[���F��F/�TC��|��;ٹ�C� = Й5I��SzN
A����j �Y��r8t��1�:�9����%�҈)����,p���0�2JR0��]����,t;g�(������E�̍�����DPVʿm�r�1im#>z"E���x<7��$�B���RҖ��j�_�ŊwD�pk���b�}��y�Ip@���:�����h�S�7�qI :�н�\j1BlH5����:���(~�~m5+S���x��!eΞ��x����!�g9�<#��G��T�-a����3���\15BR�����@���\�p�ly����z���7��\�[΋Z��~>2MؿN������f�����^��sV���ݺ���xXU�S��p�Ǎiz	H �r߹x�*6m#�����V))��Y�%V�4�o��^t�|��
게c�ʢ$RI4N���̰�U���tQB��ǅ��8����XI����W-->�Az���+ s#�`����/J��傂���`��mEs*��)p'Y���Bx�G|��܄�|�޽��S(��"��D/�`�$���d?!��K@8���$� �&���2����a�iQ4�)�?ۋ�(dmϱXI*u�Vo�7�Q��֜���B��Qʹ�_ L̤?{"�VP��Au����Pm��������͙cmG&���g�q9P �e�����f�P#��ޢE�Qra�K����o�-����Ӳn�(�L����Jrg�v��b�c���k'��4�O�_��E��G�$
)�h��N��s6�X�g��%�cw��H~�u׃֎����0��<n�g�a`El>�n~c ����[���QS�b!������iL�@3���NŻ�e�!�-���rY�G�@��L��|�4��B��}�S�qz����Q�/"����?V=Yj$�8��ߔ�nX_ ��:3@QNM�-Vԗ�\���*��p���X���ල4_� EL#w�A,{�x��O��Ó��?����ډ�ppR����_�$�I�u�I�mh:)��j�8��o9M�{�W~	%7$v^CC��S_?����\��>���9�ʭ.�0��U���:�?'���D�4��	nTj5[���%�h�H�V��Ex���aT����NK��,m@M�G V�j�)�s�
��m5�6���!�Tp���o��.�{�[ qݗƞ�	����$KP;FL�,�T������K8�,�� �p[�5��<�)L*W��1�~�� ��T�_��>�f���v�+a{k�S~��}m�q��Φm����^��˯�HE6�s<#���}rK(��f�!b���%���'R���০�{��=R����@�n����^����~F:�Rs5�����+Zȱ\��F2�}�?Зv�Z��+�^3,���;$^bo�a����8�Ư��Q�Mm�sUoD9����k�Py�z^\�?�^^g�'k�;�6!�������5E�`��G!A��τ	-�0���P���
.FW5���a�9ؽbC�-�>`4��f��i�P��e�T�r��e�H�����P�,2�X̞dy��!�6Vg�rq��Ht�ѡH���a�^�y�2�'���e\�._E|�t�O�buc��Y��.r]g��
�c�v�~<>����CU��v�%�u��z�s��(R�Kub��Zo"�W0l�f��E82��Z��h��͞.U��R�~�'���&6ߺ��܁|�����y��g��Yؔ?�¬���C���g�JZ`�E�bݤ2�@��A�����
��������S�߅�������qU[�G�G��eY�?�7��z�G'}�iu�{mc������@`��]���&�?WlE%e���f 
J�Y:#�=有φw=���������.�uC�$�2�t�HTB;)QM�jh?H�-.���A�E����652�Ò�~��F՘ ���w�c	�a�T���xV�S}�3�%�n�4)�C$��7j�F@ܻ��Ώ����{JwkI�<<Tr9n��
F$��!�t����(��ə�]#��̅9� n�x���f��Cl��S���� �S4@�F��S����F��X�{��I'�'6�N�~{���RF�9�T��.�G�c��>���.#Q��-a}ܱ�Fu�����uDɿ�����
�iN`o �m!�!؁�i�O{����̴��j���7���\\�4���u���y��3�@Cű)^��\�B�\Xo�M���`&R��1՚��l�rcF��4݋(̇n�x`�C��:�[�d˾}vvM�l��Ė����ףh]U��ǥ��,��ج�f���l_d�Z�۝W���n�"���rÍ��+�+�h'XE��EI|��@���q�m���H�;&����5�r���:�/�q��I���V���U�uV�6X��ɀ��n��a�������Խ�8Z�����KC��
�%�Wv�Br��\Ț�3&���Ҝ���hK>u���?T��+ȼ��(=�%9:#b��iC���9�O��ܭ�h��8�U=H3�a�W��9�-������)h �z_��V!4T��R H�F�3Z$�j�ʾ�*���s6���o�*/ؖ����C0��QC�)�,j�~��
�t�B��e�B�Z���^o
��i�9,7��y���0<�/b��9���!&�/|"Z��e�}��(�AD���#:��uX��t���ێ$���7t^�Ot��O�p��Nl8j��})���1��'}����孅���0�.���T
z9g�&g��ʧgl;a�1�y�AL??Zmi�{��Dq?%6\�����F��U�v�"􏜨�Ɂ�̊��O,�^���v1�|�����Ln����C������*���8�����Z�B��7H��	�K)c��g�o�l��j?7�}�s�?�7Zj}��yX��B�=9$&�L����U����|@y�/	kE|g�Z��s;'�~�0q(v�?i]�Ŷ!V�R�h��.$2���
�af�6��]4-�䏵��V��P>��$B��'��\��6�h��"������ �����A6����Ŭ{����$fk%����Y�FK�h��J~�G�x�r�qED��c�(��w�/�1��E�*XO�J8d�\����t~��g{�e�b���L�/�%FCǘ*�_��E�oVa��l��ʮ�sa�l��J^OI��)#iÁ�`� !f��AۊriJ#?	JL�?Vg<y�{��@O������6{ �t�d1L��������kw;<�[j�9���%jXW��lA�"T�u�����l�4�E~��61i���?���ȕ�"ݼ�K}zQ$�B妸�cT����x�m�Gr��%�H�]0��:���� U��I��̻�<��4��T6ͮ^MI�5	}iqp��P��{{6{
%\D� ������^��v�����+H95���]K��PmqA���o��K��r�V%�������;r��'�o#m�n�a�Rs��x�ڽluJ����A�i�e�&M�MCr<�����.�K���|*��X���ढ़=t�H7߻3@�ҥ�K+�b�f�����i�w�ql�5!DD��d!u�������L?骚�zi "��G|��z�*���m��}+(o�J�E]���{�������s	w������^�%�o�(F�m
w#o�؀���/����ue���*LӲ��i�ߞ�Z����-��<��⟻+�N��JhI��Z�P3���<?KH8b13K�hF����ƌ�
���t��W�����ԑ\�O)��l���Z�
M"�׿� �s.������z!So5�[���n�E��h�W�)�Q#��k��p5�-�μ�#JFN,�25�f�۶G!�v��3�����_�jzbQ���W����ޣ�óE,���U��
7㓞V̆���%��]�͝	�����jxP�5ʈ���_X��vFJ���7L��kLq��^q>Q�s3�a�uwkr����,�7�T5|��"��/�~�W�|���ե��a�2p��"�?��n�AW\U~�D�s���l|�������+E=칎�Kjd��Zh|&��V��b��V`wӻN��u����ڞ�/
R�y����=��#6�7Y��9v�v��޽}��K��~9���󻱽��j�|��:؏� �u�>�%���Fr����i>rm8y���r�j�XK� �j������>)�����ݲ_Իd-w�V�}7�Rui�fm��-����Y��/J���r3%���q�:|�D�B�;�1�W��f�S�+DDP��h������:m-�f����˗a��3�;�&�@�g����3RqS���x�$�)]�/PA�k����e�����-�Sꢅ�xP&Ԅ����KluB�{i���Մ0j�nMv	M�&T�3ZZ�TU��������=�>I��`M���(r[:��e��.�����a9��q�W%�DWS_Ĥp**ǻ9*�gW��WҰ>S���S�|5T��?��ھX~����>J��y�
��t�	Y�z���8��7Q���Q"E<����	ӥ�S����c�ŷ6��ѷ����l&l���9%qvSc�N6�Ow|�X_2.6�x��n$�L���_$:���U��\~�n�j����d,��6].�
�9^q�).�ZW�j�VR|."Ȩ��S�R�,h��-ۅzߋe
g����xТ�"T��+YP޾��Nn?��j��L뙕Qѽ��n+'����sM{��M����Ax���(�r��i�~ƨ�+���J�l��z�]-3\�H����7��Y/g����'j���������kSJ_[�=ɒ�m�%�f��Ec�����9�<��f���}?H�������Cpק���J�U��m�B���2y�IÚG�Wx�Y��^qj�csV�� p�9l�hp�v�n����R��Z ���fUf��Oy	��$�}z�^f\3��o}��YɅ%x���C���~#9�0�Yl�>�{�)�RdK��uHw�Y��O�?�bnc�l�GT���{��|�]���|��V3����Q�sj3M� �U^�F|���>��v(�����a�uɜ������p y��c��u����H�����n��"s#Ȗ�깊���߸�v��Ӧ��zke@
J�Iz.7VX���-��֒���V�\����>�1��d+�X�T�/b��0! 9��*'�s������� e�Bp'�.�P��h4�eh�� ʬ����c���|�D[�����+�}�U�(W�����K�۳�b�Ԓ����Q'��=LB:ɵr�ʇX�Z�T{���!C�%�l�ڋ�*Ұ�Xq�X!`Y�g-�!Ky�l�R( �(n�\ޖ���V;F^*wq�D��Y�M ��&�_�hjУ�l�Y�X�ʊ�<M��C�b�Y�s�|��?j�*R]eF�1�A��'������h���]5��o��14��\_���*���Y��w�L��}O��W��ΊB(k(Ǧ���F�-��m�AI�M�8�� �	1���sW:��T8cz�d��pU�&�c�#�D�],-���\�gp���5N����@���Lva����J�PSռ���ܒ?��U�x<rAµj���Nױ|.wk6ZB��ﾛ�C��*8�]tX�i׭��f\��B����F���!�� �K�Lײ�������V�;�
��lV�OcH]��MH�%EBL�����/�>}��ޒ�1�ě[�v�,,qL��ء'e��u i9�2e��1ұ��:Kd�f>m�����X��&���%�k���� c�m���؛<�γj�#�(���eƊ��f�{X��(��-*���ꭀ(�|��Vu߼����vmy7H���t�h��H�𵺟���Py��b�z��vnwDr2�}��ۺ���s[�yY���4�C˦u瑭u�$��BU�$[�iB���f��(�z�~��5��F���s�<��+��P��9���I��7f��J���=Z�cѫD~��g��en��I���4�����;ߥv�ڵ!������\��V��b& .UqQL��p�j��qܡ�u�X�\/ i�[����ݼ�kL���{m��V��ߏC�t��xh�o*��~{'.L\C���"���h�G���H��E�+��,1 �B�ϸ��f>���[��ħ(]��W�[�b�#�T����5�
��k[�%���\=�mp����)|�A)�d|KN��eɒ�K��e��\�i%����B����������9�g�a&�L-3Am� |Da{*x��둨�2��#׻چM"L���^�E���;��KS������.�q7j����Ӿf��墸9�v��Qx�I�������˻�-��j�� ０E��iO�*1��iJu��PB��?֗)�^fբ��o��o��;� ��e������c�TuӦ���7G��~t	�z��>*��D�{����{�;Ḡh��J��m'l���gm[3*8i�౴b�����Մ��a���f��;�����k�
{���fb��>ȡ䴫2�\"~�h�H�N�Y��ؿ��Q�2�?z���1�����e��$��t���4�#�4
>Je�-S��utrǨ��������\�d*0����a���( ҽ�76����4���j��]��fe���?β��[�E�s�� ��S-X���r'���D9ט�`�["�|�t�8)n��m��6z�>E���}(čX�yv��_˨Xs��Ys����z]]^x��w�{*��Q�ݛ��T'g@�a�v��s!*]���5������9-�NL�Qҧ�@�7�k�CR�h�vlsa�֞�j���4�0?,�9�P�7���ծ�Uz5���0�w���;6��q������8�������m�����;k�p��r�s��4�i���o������Z<]BЯ���Y�S출R`돧���H��m���%`[����<��-�?Z���J����Kة�W���I����f��[����A?a�o���,�O�j(b�2�p$;�e�v !W�|�G��x��y���/l{G�0������9���^UP�g�Z~�H�b]�G�BPS�����6[R?F��ߍt����@?\�<��!�����Q��6�I2Dl��0��ۘ��Xm�Py�~!�3��N>N����θ�=�h���I�z��ZU�T�y�yUBQ��A�*�m�{�� ��*Ld�:�!ϓ��͛�c�|�x# 5X���R��ӆ�������Q*�Ϯ���?37C+Xh��9w���uBP��jy�^]�ƺCke��i�us��>̵81^�ʁ*t2f�j;�+���J�����򠮠{k��k��F�Jܹ�?�Պi8�{}��l���ԋ��);����s��|�����:���/�Vo�ūȬ���6��n*A�w�xľ@D��'r�<+*wr0���)	�t8�=�f�%#��0X^qǤ3��}g��T�6x��Ķ��$ӭ���US�o��\��὏aj���SY�FWP�;�1��q�� �d����U�)�1��谫����e�C�%ߧ������=����a�uЅn_0혯Rp������3�ꆇz�x.����6���P�x���8�����Y��De�P����C�p���z���=����_{�i��έ�����?S���z��틴n��m.�������C�Ų�_C�HaJ��խf�����޺L)ףD�4'j��`I'&���M��d�b`y�e� ���/\2����cOq�W)���v�b�Gk�`�Gu��՘M��[��͇��N��I�2�i>�H�?P��49�e��%���D�\�Foޕ�������m�ݿ�C�v8ߢ� 9�Aj�kJ��������ol]g������R���Ķ�"�bk����g ��d���j�f#��U
�/�*k-�/�֭m����X��J��ƭ�s�x�P��(u�������]l���$q�$s`+�W�ߙ�����J�W�����l�z�D�����?ѿ'__��!#�VC��S�O�	�zk<y�JUsҤ����b0�;�'���Ε
f
������Z.7�����{ A1ɖ2zwөL鞮��F�{1�m6��E�-���j[s���N�g��ٔ&��b�/�uM�*nI,@%zÔ�F/��H��1��+���EA�\�+�2�J�"�j�
4R58ŝ�kԎ��k�m��E@�ٗi;��m�΂P��Y���)6��,�YY��>��^:�I���cbU^�����+�v �X�FKk
j�[_5���n6�W�!c=�� �����R��V�#\P������B���{b����b�Ωm�.�L�.9y�7��<���<`�B����.�6}��`E_R�o�cw�k�tNm�-?���?%����v?�Vy[����F�XY��r_I���i�@w�։��q� ��FG��������M�#��fS��4�����9�ڀ썟Y�����^.�W�1"�V*���3~��8a�Vz|���Ƥ;E��y����(�J��J�qA	��W�i��n�K�hH���Z�^f8O��ytѾ�j�Nw���޸ȕ <7�v�{�Qb��%\JfQ��n�,��|�؆c-�*T}���h��|�g�7ԭ��5�|�����s߷��^6�h%4�j����'o���?�����m�[�O�0C��7ݾ��ܦo���l���=SE=��'����:�ԭ~��>xS޻��-|���R�i�u���8c�f,�6��$�%����(Zs[���+�lP�Xs�����2����zU����=��N�~�m.��O�Iy |<�\�h�cކ���t����5b�)�N����o7�v�||��ud9��i �BZ�^�>k0�
�ZXo�C�9u��r��1s͂^�L��:Z���b�x�}�V�c��8�����m7�3S���h+����R��ob�Ul����Ҷ��:�\���D���0���v���z����#���i�k�
�[���j����]�}M/��q��˿W�JB�Z���,H��r���3��+����'���KVJ�f� �C��D�wv	'��S�N�����=�s��9)�Vr��.�@i�N��������Fg��jƿ9k7�Ƚ�u=����5C}t���^L�n�����ǧ��w�0ڶ��_�i�y�;��<�sg3�|��D��]Hq�T�o�G:)Ȋ&��A�""�̕���G��#7p柩�n���p�[C���h{ۿ������
�-�{���M�+[�u�Z����
ʦ'��w�-�+~�~t΂�i�id�q���zƁ�8�����j*+v�
sk���M�WbSz�]^��BEt�c�����$��=~�\��Fb�ݰIs�W�(�ď��v']+������u�v���y� 6C��e.ܞê% ^��9Ǒ|��r��f�i����*/���m��LjHЍ��t)+��S��O�Qt��G��Y�o)���D1�;�� n/[��w���cF����0����Vܑ�<�q���;�۝Wb���H�z�#q`x�(�$vV�ZPWmϹ��LrM���Y,�����L=mG�L�`�-�_V�f��b���I�&7��c�fLp���v(�8�gc>0V��)�!�8��b}#!=�6�y��i�a`
ⓍZ��uEPvH���<����@�^���k�)^yi��h$�?���̨�N��h8�S
Zݷn�5��_^�ީ*(�y�L|��5_�2��<Y�c��d�.��{����w��ƶ|���$
Y@hE�� �>��6�,�e̸�'� I��[�
��m'&��0(�!�'����Q�Bhr�i}y�χ��������r�}]0�~�U��lh����!��o5�3�E隽T �GKMɹ��k7?ѥ���5�u�0�#�������R���B�*���R�?׎�˳;��?_S���惖UP��n�0�8���n���Eg�:�P5!�?`g���������鞇�t�Ʒ�9�����}~���vf��/6D��>|��זC����H���?#`ZY4�JK�vA�����7�;���1�G��,4f�!�å����g���.��S���z��w'$���_����y�/��1��74q��s[tLw 9��Y-�1���"�x緛����Q+v��o��U|K�'�^c?Y,H����?<ϯ�T
��[(��w���`0�E�r�O�ٶ[�[��-�w�,i�a
޾�F�y���LR�r�_��/�6�YK��f!`��c�J�l��=�S��23�o���t�?+��E	�\��g�����\1�({43Ѥ���Wp�ҐM�����̃���֕��w�އ�����\'3F�5\���@����f���e<����4��	����&�T�O@}1�,��.��H1]Q�u�T�;�(�eɾ�>鱩�P'������Q��2�d�yv^�9.�V�g	�O�����+Zk��$��>y���O}��gqqG.�p�4�4�fK�����6?�c=V�3`��ۯ�3s���u�����w�E�l�`r��ł0@�~C����l��n3�L`�Y�}��@s�7�~:ZS0M��4s�WƸm��S��u�r�ݚ�f��HLE%�R{X�qC���(��wA����Y!/��/�t�r��Ҕ+�^I�;z�dx�F�fGS��0��U}4����UI�3����f�P_c��!����p��j��e��e@t�[��z�?h˝�����������ʢ�ZëU��UG4�oo:?U/l-s�}pAQ8�hI�j�^�'��a���9[+���7�������qt&�^�80�R{��WA1�AЄ2ʣ�����X]&���g�I��;�ݿ���6_�&�Z�xT�w�%�i.c�o���1b�`Q�ڞ���<،́_T������)��s5���x�d��'��v��T���&ʉˬ��44E�"Z�j>�U�Mc#4JL�v��k���s�Q##2{g�G����\WU��Z̏�	�~r9t��8zprS��MrDe8�C����`Ȟ�>8��+��m�j�[cY�Q�����B��-:���땺�m�9�Ķ��ڱiF��f	�}��k�ր!q���~rBم�����{](�B`fiR�.�������}aa&��tz�����k#{���#s�x��c�yF{��	���E�Vې+7(�������SԊ���G�`�Ƽ7mPI��&�x�Z�)�Z�$�Ժߜ��F��I�T$�9Α��P���!4��d����$���<�ye�XǍ�����sK����J���Cl�V�@�{4`5Ԥq���A��Cֶ��X{��s���^P_�Y}q�ڳ�?*��W��㙙�
��j�m��U�y�p�ػ�s=�:U���;OvǔW��c�p`��i���a*�6���Y���1�ɣ1�V%�OڞܟG�ec/���a��5[l$� �e��l>��7�៸��\����׽}�p�*�@�^o�cc��n��l���g#��\V��f�e��L}&�I�3F]�TFSW��G��9qe~��tU�M�-A���Syk���j�ҩk�aq�ZY-Qג]���i�����m���OJ�-�%�7wI��h�6�	}O��>�Z��\�#���ظ��d)ť��8
�F:�Zd���b���̧JcEE6��ݣ3�I\��!�������������K��9�m��"��x|�g*�rw��.\�����̈x���i�A�D ��n�����EQZWq�@
�5�.�/X*R��P�dD��ET��d!�$I�؎D��;��ڡ;	cV���x��`�2s/E*{v�lS�]���k�����~��#���?�����u�ARM�?����帍�26���1_�3���i(B����S
!�EG��\z���-.*q�`���������_wk{��:ڳ�^��# �8>'�t%�~��つ�Gs��VH�*�A#M���MȧUB>T�H�Q����%��3�C���]����2 �XQ��'~���̙�($�����ss�$�=b��m�� �b;��7,���~���}�;Z�n��|/QB�F�M4h��$�C2`�_�!6l�f2�����?����.~�#C�a��(��rT"4B1�����nbhy�&�l���H�����k�E��\�l�it���k�e�?��i.�v(�R����:�:�z� O�-�niu��r6 v�%@+�yU��wg>���ʔ�+l�<�V6_�?����Ș_��mq& O����6{�菋E)ާ��2��v~�2�?}��`"ݹM���llĕ�_����T�
��D;�����M6�"��O��@�xr�>��b�*��������J����ϴ�/F;���߀w��8T�:�5���~X�Fx��c��x�f�3�$��@����f�������&�j��� �)q�شEnlϝ�׻�W��7��K=�K��d��bֺ'.vJ�L��t��;���rDl		����ӫ��ҕ�"�O$����3G>�� R[�y��F8����]�˒��=5���-����9���C������$-|�`�5�����'�����g+B�X�ߠ���ԝ]�o�� �ͧ%!�=�[W��ryD1b�|H�/[d��֠FE�������u ���+�y,c^O�c���?(cƍ�$��}�U-�W�x���%t�R�%c$	������
�C��rz��#����CÆ�҄[��CU�(���
.��u���%��"���~�����-�"cl&i,)1A��������������^�7ŷ#*���.��Gj��Xj,����̟[)Z�7��eKK�����'KI�h啅k�`�)
WTqh�!��P��|y��r�\A��h�$�w�Q�����Nv��;����h�^S��Í��̸7X���n�Mq�G�����RNe��jÐ#�
ʹ2:g�W���g���l6��'��*d�zJ�/���'�P+�?0���a�Ѩ��S�y�㈸�h�I��\�le����%�>;�܅�#�&5>����QT���0��rЯc���<ȏ=��'0-�B�6�av(�����^%�h�Gg�p+V�ĉx�/t�ԗRG�o� £���Z.]�����*	n�#�u�7ġ2��Я���,�_D�HvE-�n�
4��ku�2lL����Hd�Z��ϫ�> @w��%��7��d�˔�Əƾ>�ٶ�"�'W��JqL�I��wi �x�1*��޻2 ��o!����򿧕�s`\��<sn�O=ߦ����g��L�9ݙ��Pm@@P�E������f�t-	S��g<]�^�����y�k��$7-@܉j�9��z�қ���ӏ��T"�������Vݤ|�l��c̲�5�'tɥ׀���bW�F|��7$*1z}@��i��po�������6��1Tbc�{�d�@�G�q
E�n�$�m��o�����5�+*l��@�ES5��㒀B×��0�".?)n�Y �T���&�op�u,!R'q��V�(��*���7~�J����1Fk��ۃ��Bw��n68�m3X���<����ޅ��5���fQ���9�jV���hLg�^k	�(�&��7�kU�mV�k�E�>�fB0�/�>��YYK�u�}�%��2J哌��bijs��s<kl��Ǣ�y�y��T��e½͵Ւ��:]���l��S�����ڡ��� "�1K�֎Yi�g��/��=4hJ� \�%�c�TR����s�����cԅ@t"<�r��=S\7Lk>�P��S?�g�#r��\Ur"��f�c�e� Q)�:��e�Ð7	Sz;��CY���D�`�f��jJb��N� ���@N!��fmXm� 6l��}g���}^CKƻ�^�����z���	��q���lT�F�����Laݚ2l2��T�y�kb̈́I9d��r�͕���>C�^jWD��Ga9����a�DV�d��5������ѐH�M����EB�ŧ[�d[�RM&�o������F��ڢ�o���Q��M4�����8��4�����v������O~UX/S��~L!~^��2�+r�{8��1tk��Sq)���5��<�\.­���`˄*�Ֆ����m�v����?��v����|�3c��?�B�#����7x���!u���3I�j�3i�����y��a�nc�P�~�.{��|�����փA	� ��� �@�Rɻ����@4����Q9�#z��B�ۼ�;>_�x,j���dF"�陓�k[��Y�������R�GL��$���Cۉi�C���
��'��5����V� <�sv��`���^� �w2�����X\g=5e�0�5b��J���6淪��{8&��mFۼ�����]X,W+Ǧ��UL�s��{�~��4|����k�PF�R
3Ů�jȃ�q��|W=��+���6L����4%M"��|�+����;�(�G����q�*����휲`���ݮz|�̖�w(�u5O�,�Zj%L5c��;��gW'��oR#V
�0Ό��y����#v9,R9���M/5Ĭ/kv�a�F��n�֍�˜v��'��u�.~<���+?�gcJ������<Cw�7B�O|+Amg�X͑�P}�p��u�O 	))9u^���Ń��T%X)��<}���G�30|/�fl��O��n��k���ӓ�ԓw]�^�fĩ7�5������j���a���Zt�kh�o�"P�� Q?����J[f�q���� ��{^�U�'7��*���>>J�G n7X��W?S�.��V1[l�!}�w4�iD�2o�xӔ��-����i�tQ�]��7��JB�����_;�
��돀\Q	?4ײ�p�}r����#$L��u��w� �V[zX�T��+�H`^�2U�9�{V�MBG�Ps�� >p��th�6W�V%�gj�%�]���*�U�D^X�� ���~1�������]���ҩm夶��7��<k�5'����(#5�Å�L;!d9�|���w��ߘ�8u]T��駂����&��B?ٕUӢ�2G�
���M+��H�����nɘE���]O�f�\���W"QF/�	�S'��3o/��f?�h:�枒� <��V؇��f��][��㬎����Ua ��$���|O4�:��ɖ}�ؑ"����z�g�Rt�����#�ن��޽f!�Mu�T;���b#�2Ƌ�_M�����1 wuc��0��~�\]�����x�zuI�n�UC�܋��H;��C2(s� aȠ���'Y�!���4Y��'��W���D~��dq��w/oM���ۄ�j��h+X���	����>��8y�.�~䴔.�_��3��X�H�Ը�N^,Us���O0�H�>�Q��k��6�k:��E���'�$8g����!H
��~�4ȭAw;E���0������3�֝�4:6=�*�"0�(_+�_m�i����p 柵�o�G�:��E��4ԐG�d�b���H>bv���uꁓE-q������ ���G����TF���D�����f}�fY���&{=F��E���VŶ@���9�(����a�!�#}�|���������X��j����+H���U��V:}Uh~�Wi����5�-��N�be��}U?��C��K�8B;m�V�N���NL9@�5ٓ�6�)V����X�P��}���Ӽ?��ʪ��;pγhT�D,� �"5��K�{F����Л'"��%�r�ł=�R s5���,1��	'6��w�_D��K�
P��wO���������y�Bd!0ZǾ��I%Ԕ,����2H�Zj�FS%����ކG��=��3J\�b�}���X��-���=�`�%=F�o�'�	�����'��;�̯p���zDj�|]�T�fZ��Af�Mل��k���	�?���s����p�M8���UTTT$��$Ǧ��TJj��t�CD@�%)���1Jr��k��؈�����o8��u��ypL�O��dg �X�Z����kM�[Z�l�?}SL<Д�|9TR��塁q�iZ^c��ܝ7��2q�l�iFO����]����f.�>��cq!��N���#,O��^�3�nY���MlYq!e̏��a~�5�cC�P��_,�v ���R�I[�_7q��J��۴pw-��� �U�j�{���X'�>�~�k����*�m2�ggh|��i�5�fإT�u�GMw�����d$�N����qw���>	�Ep�
��U��������Q7��<M��4�;�`�3�-Mu��5�M,yῳ-͋�qנ�,)���XS�౎'#��[]��աF��UR�y�X��|K� w�)���$��H�n>��#AC�+]�N��K�5��&����-�.�P3?�ͣ�<����C�;���Z��a�,6ej��q
��y���55�~(M;�-�l��Iq��>�F�gw�#n`��-���RTm�Z��G�X�m���?	�e��G=���S/���O�f��3{4-i�w;O!�s��Z�[�#��W�x��+F��k���6w9�w�󤚦 e�uPd�<�/���>-�H^���R�@���\�U�«���Na%tl���]@a<��+KVݑF�R�B;P�@W>�n׸�Ny�B7��:t����@
f4#>k��C��b&���^ e��~(%�Au�9Qm�[vgD����6ղ�U��v.���	h�!��A]��G�sN����Ue�u8##~�B��3�B	��W)�$�-��L�u���	�i�ߔ�9ˊ�=R<A:x�:� ��w��8����\[i����PH�.�w�	L'�;}�VC���a-�-�98]�IX>�����X�k����%�H`{�P��I; ��4��3F���ק6P��A��7#��n�+)5�wVc6FeF�9JiAw4��p�E�Ms��j3Sz2N~�H�oR�c*�p����o�6��Z �Fe�4�@U[��k�Z#�Wz�@��	�讨/�n���e��꣒u��ʽ�?�c$��
�zE�E)�y⥈�~�8�!������ �lsw9��d~�"�?�)2h�S���+�%Yi�V���y���52�B}����'�*���%�*������m��o?=����2�/�f���-tP�ז�X.i:���L-�M`_Ll,y}�o*i�O�p��������5� K�l���^�c`I*�(W�SAb��ܣ)�����= �Y�,�)]���w����U>w$غr�66���T5���^�[���
�3TR�#Zغ��q��>��@w�b�8��p��CAN>�+� �����h$=�����Ĭv'�|g @����T���rš�Ӹ2���8#�t�`eB���]D����V��x��
��M����Z�ٿ>&�_�f:�(�x0{t�+���s�N�D��ykT���*3�|�g�}W��&�A�O6K��X&�:m�����/����oY�Wre��I�W�b�'#~�ĵk�  �&[�!��?!v8t�e;"���Ӵ�s`= p���|�[n�Km7?�vi&�(5ҦԶ��zhљ��Ϋ���m*���e�&U�"�dq>x��jl�8N�{�:2^����L��3n�E���/,��)��r#E��N�e�4��R�q�W��m�V'�Y������ES̆�m/G<���A,��T�������/�CI��p.Z���}���|~�����Ob�����o3��0�`2���4X�Ȕ���j�"H�w+������ G}7��-��#E���.4v���`����w���:�R��'TU��T ǝĢ���W�\b����@=v2�S�Y,�ns��#,�a�����U�,ғ�||^ł)���ʎ'�R�I-R�1ޡ^�G�忝���:.-L9�h1�|�TI=�/�ӛ1�J[�Ѵ�ތ��O�%�-��\��b"����W��܍��=X{���1�!���VvRqu.��V: � ���f��~���Ìn2���o��N��6�_�
��b�e?k_�����ؖ{Q�2~K�[e�]���!�o�O �~�V����̎Q� D~�I ��r��V�'�=).�;��'X�R|����!�R���4���ؼ.Zqᤸ�<XUEϘ�kl%�c^߫%)��.+�|C�O ;�R���.���~;i_��:��S(���B`l�2\O�?�D��o��9�>!N�5}~b;:�а��F��-�9�^H�5��W���T�[�)t�˹8��hY�3���R������bؗ�2Ц�7�h� k)q$I��{l�==���K�5�3j��'���&�t����y�"�<��fw4\)4���/0�=F�Ć؛h|�{)��\��+�̗�������I�}��=:I���w�9;qϟ֫��eP:r���kW�o����o��#�� �.e�����4��Z�;w@p���mc4Z?~����<N�����߳�^��f!�����~v�	�ٙDl��z�y��MP���s]|�n�7!R��4Z��i\�0�I����U-]������w�6Gya16�d�ر�܁��;�_��B���_�'5ۜ��ڜ����]Y/���cvzY�������\]r��=.>����r{n5�(q���jc��_;�c? 3�c��e����5�Q�I�d���>r�l|%���V��e�G_U�Ms��|�t����"�\ʎ:�T�U����+u�Of��V)ّ6��	�Ε�J�}Њ����`Hg>?c�}���x!�\n�5`��_�͎��t��X��֏�X����G��jlӺu:(c_��E�1o���ۊ���|y3B�\*�9IDߵ�����Z���wݳ�vq�Ǻ�ܲ�~��*�'7�[*��u+87�&�ln������9���(�k��;�s���˒N��x[������W�C�c�L��Ƅ����k�B��{m=�7N&�Nn���:(>�����+��k�^��=!���o�����l�Z�����lp��d�&Y�+�k��|��dMIƆyU��s��(Oi��x�K˂����Ÿ��j=������[�I��);=G���S�JS2�'�^�y��*�F��!D2i�:�F6��V�L
w�T�Və�ѳ�O��6-�D�Wt_�ήO ��{��[
��l�M4��b��w���<YQ'a�`����8�Z�D�����Ed���w��g�ɯ�ƕ���U�)��'�����w�_CŖx8�P�Ƨ�ȕ�yV��;Zuz����y�Ъ�gJxm�����䑳?˜�HY��ݾ�{V�����q#��%v��J��o�ce�H�`��W�{�kŇ�i���V�ﵪ��׫؆/�nn��q�"t<Ik���Q�]�0>3�m�������3toY��7�jr@�b�{�sJʅfVЋ�k��X���׾�V/`����[��5�w�*�@����.ߢ��ݐ�v�.7\e�:|�n���L>���}���Ϳ.u�� �ť˹��+q�A�0�ߚ��p�M�XIB��0)	@�Y(�#U�uk��)�mkш"Y��i�G-�rTO���@@�Y������t�KaV��74o����q��tH��e߹�$��6-�����^���n�N	D�?t#�h)�r�7���_�_©����W�G�;Ŏp��q���*,�[���k�c�8����9��=�#��J��J�R{��x�w��[H�x4�{Ba]rkk6���[�*(otU9͖�v�a��N��z/�-��䆳VHꊅ�����qCbiE����J���F�Օ�\���l���7)���t�x�2��]*�t-C�Y'����5\ʴ�v^(إӇ��徝w��8I@N��x�obA���?��r�"�9�%x���ʫ���?K1���TT��y��]W�6]�Zy����dZ�3>{��8�S�(�����w�\SY+E��>:S���^�A�a*�\ćg�ǯ
�^����X��GnjD�bwd��xyC��Jp	��-�s�9���dH���� ��|��Q��D-�I
fA�+���l�3��m�[�t�(�UN���Wւro;Q�,;����*�qc���Ԧw.j�u�D��E�ޙ� "q�P@:�a�|��O�Q<�!*�3�}����J��2t��hy�5�Q�u[�&.=�,O3��Jk���7K���
z��/�>uFy����uҨ�������s�(��y� �o�.�������@̏"����s�s�����g�ǵ4�+ �υZm��T��ΠLds)�?ӏ�7������͟��;����YR���i���mB�:[,��%��\�������Z���_S�_9:_�E���uĔ�l��x��!�ca��{!�J"ԍ��s��V��s�W�Ɩ�^�r��`��G�s:;Ʈ��Ζ�4��7h�u����x �#��X�3���{=f�a�S���"q��8d�C4�N��lW +�����z)/��>��z�H�R�m�A��ڒ�?[���|�s2�s�c�M�0
��^X/ݚ�>����r�J㸗��)3�ē6_%f�y�o������צ��mv좜��b�F�?�k>!�Kj��hpLAq�A�s�]�3��=��V&���#&��UmX^X�����\���l6����/=kꧻ�~!9��ģ�u�G�D���$o�z��P�"al䊶)?�zǟ�9�u�sV��u����-���{�o� ��7��Ǧ��ݼ��#���f���.�<_�J�m�Hz�aḞPK��Oj�<_���l�K ��wb�gd�?+R[�7/}��Er�[�YI��˾�ZxWva�p���^!�w3�̲\F6p�K\h�2C�ڥ��
����'�u���r|<@��	+Bu��I͏d�u���K~�����R�$�8�����
qh��>��?�;�ص�i�\ă}��̽v�I�6�����j��Z���x'sh�|�����e&%���]�����ٿ�����S�@>Wm����[�G/j��~b�L|�w����I��/��	�xv��s�m�S��ǀt���ѱ�����_�យz��c�-	���Dxx��/Y�}�)��t1�'��X}TIs��v�� ���6��S(�ܙ�������B��9�q���k�D���1I���+/"����i�����.���&E��7H�]�S)�����c�u�Z8�|�z��;'t\�۲����9J}���9����ZΫ%h���E6_�>Fz���L�b�j,/�S�����r�?}�>I��Z����Q_3,+c	�s�?�h������oX����]�RӖ��#�hsxLY/�����t�Q��ng���]�#�X��.7����m�X\�SV�tQ}O��~��g����4�+$Sq�?��m��6H�e ��  ��������~�80�e���-�h�r�"�s���7��{� �^�BЍqZ"��Qa��Š-j�+��o�*��Y�g"b�eѿN��PT�}���o�n�p|�a��A��VA̱��FU���o��c���N�6���BV�є�ENhF����7�4�Uԑ��Ɠ���������AH��Fx�����ߏ�E��2��}�D9W���V5E/�����r��Q[�6|������3-�u*4�L{\�������b��Iw~����jÃ
�,}��c6@΢@�a���}�'p-��ly	\%�?,�#v�K��ws�}�J�$E���A�/�82�R�5�?�Z9kE�מ�s�훓!�7}��/mM��Em�:x�=�z�+h^d~%2�)<i�
F�>��k�4Q�zq����'^��t��L>��(YѢ�<����8�b��5����\��V~�P��qLh�u�����!��'U��չ����,G���-���F)�]ߘ&��"�l"g�b{E��v,�ƪ��`K90�b�gDG�
�{\��zJ��F)�Ie�b�-#MA'�~�#���������mO����
�n?��J��n9(�Е�+W�
��KZuVM�Wp�y�%�/�������ܾ�m��~��{�\T�٧+j���pr�Z�Y��UMNj(�Se��`V�V��|�U}�U�V�C��V�£���	s���\�����A;7O���w^��uJ�}��-^lC���Sg�����oK{�	��5Y�Wr9K�HR��9�OA�RH/z�6I�C�Q%QB�˷) FE�lF�AQ���"�H?���u��<�����[� }�ˎx���d��v�\��äBmѬ���Z�&�s�pxk� ��RS���]�t�*�O���5ᣭ nG�5�j��XT���^�d�h�ۃ���%?�L�њ�_;��]E�Ңj�?f��6� �J����n�2�%�	����m����d�T3���]G�K�3Gh.7���m����3�^��w�|���1�����Xo�m9����#����	3	Tӏ:�.��M[{n�k�wIz�f(����c߇#�LQ�������L�0�ε;A;�� {�����|���Yq�7����UX��������-2l)��3"�u�O�,��@��o��a*���<���fm�o�᪅e�V��n��w-_���T����.8$쵘M�n�;8]��w��n�8І�Ը���߅����/,d.�����Yg�؜�I7��ǳ�q�5���sוg�B$ &&�˶%ݭ�9Qx�%�����KqiH�/��<��R4���M�x���AZD	����hs��_�D��˵��"��\�����������W�1��:��Y6��~%�QD�Ë�@/P)�a��I��R��F�1ƞymlP fn��vCI(;X��F�8fwW��̽wa�Ux` �8e]��?S�aaw=����eg�X�*y�_t�fm�� �"Y��1t�3&OD.Gz��	v�J�%�~qf��z��Cs&{�����M=�@��`��T��{�Zh v�0:�W�����Ex\9�������y�p�9��%���=]!�bU2p��s(e�Z�	#s~n!e�x��*\Dɢ�Tb?lv��F�	��{:�-Hm�x?k�QC'�E��0ך��!�������_��T�أ�����g{&������"s9�vU���R����@����n�X��c�E�4�/)�'�[��(#Y���߿!_.!m���7Nk^=����ߩPx�'8o.dahV��0X����o�EW��7Ac{�}\g���J����C��$�X�w�;!�2rY�3�A
QG�nvs�k���#��ê�N@�<�#&)�\8;Y�h>�����⛁�g����=�!z��Ԧ��hN�Ҍ�Ih��e��=�[��bp��D��vm��ѧGS5�k�����kC�j��ٛ��曘c�@&���tt�b����{�1�{
_$��Z�8QK
�9��ఇ�Wk4�sA��9�g�`�m���Y��ag�RP��T��;�Z���U�@~�У�=@\��{�%S_z�ja9�3݇��&�3��)�_"R���O��얽�cZ�Zϙ.�a�������@�����������˥�gt�v�<b~K߯m/Rz&��Gx��ׯ��k�{.fCkMOh@s�2�S���@� �(��N=�Q����`�n�X��/>Ǉj1ŶaQ~kw�mQ�`����*�{�_��̵�ϣ�(.}��ξ�$�%C{}v�6��p$�LR�ve����\��<����'�����/$����ہ��j	_�n�QL�0�J��Ҝ��k���R�9�@����PrP�'	8���M�C'�IM��/�<��S�ln�$��|�q�C��������ױ�CGX�dю8c�n�3��ܱ��K����?n@/�
�}9@fԔl�
��ځU��8+�l�a�G�{����8Uy����!���U�ŊᨘyՆ�����?�.B�[�ҋ���G?D�����o*�B�0�[wvM�qR	�ų$n9 ��K�_��&�����<Z_7UP�{Pn�a�����7tH,�>�Y~��6S ��h��'�iTjG�A����A˦D� +!�6��EC1�3-a�</��ݜ����p���8٫G:�-,f�[0L'�a����忧��N@��,��a@�Ub��LuSSO0�Y-]�;�qC2{�#HIc�Vj$��C�C����v=Ő��w�A�GJQ^ti)�-�������k �Z�_��JRgB����5Xt�*]���j��	�.cL<]�o�|�I#u��P�`9��(�0�����S&����;=�DQ��>Jw_�}���7��*$�Ae7X�uB�ubk�M�(3Z#�'6�^[�w5vК7t��@Lޞ�Цì��	&��{�]�X�tF�E�[w[D���d� s���e�����^�x2���ng|����;�����qbWo�I��~��I��+@޿��7p-qZ�x����ES| ��z��U�$�m��M,UQ�-�����Ƞ�OD�+TBe-���V��V���q�ﱥ�����1�,����C���|���LS2�o"Ɔ�/Q����}$�#�Ƌ�2����Z�"|�����wL��}zY��&�tWe��&�?�J���A�ª)����ޚ�̺�2���β[$���.�w'�M��x�
f.|AXL�@h���8��a�'�s�0��m�SA����|��#ڮ�Z	���l,��5�C�S��̗�D�\�1�$�9Pڋ$�#�K�&�T"J�KA��RI��L.P�J����@�4���:����*�r��&�i�r�����]7�H�F��Ъ^��~Pk��A�m.�����B���l|/e���H�ԙ˚�R��y"}p�ΔN�����}v��M2c�*tvV3��Rjz�jU9��@�lr*�?a�h[�g�Z��D�C :F�VC7�䶳�2��3=E=t��oa�\*�)i�u<�
_�,E���ʱo�^���'w�#��Aӟ��aC݋��si�.%�])_���֥����:��W����2o'�G�*X���.��%'cJ@%t1�-�*{s��	��o4#xݦ�������܁�O<���x6��A�O|�����nR	s��-��6S<$�S,�����V��c�(x"��Bi:-=��3�H����|c�E����`����UJ��\�ܝ��(�ێ��� 8~��il���K��@��θ
z?�6K>%���j*.�I&��'�l˃GaN�(�s����7�H�C��7|{�+�`2��C���̊'�]��Y�I��̺�փ�o������W\��Msב��u�(�:4k�>�f��MN�}Ԡ�x/�Y���[�ĥӧ���oc?i�˦~�i!�x4��u�pm���t�bX�չȲ�״��K,����
��ā���-z_,�t�u�Ly�Qu�����]��<0�owm`}Ɨ��_`�"̽� q�B��[7����(x�u��#�'U�~x��s��O��c��	W��S9����>סHG���\_^Gs�c�(�]�q��[�^��H3$mXT<E�ک�>)�9���� �o�U�K���G��w�<�C��C�+��17]K/xo�H�cIyu�Oʸ��u�@�?��+O�uu�Q��׷�i�>+���J}��z�xk� ���ZI�%o�q �aŖ��	7HU�Sl�␬�J+v)����<i� �OW�S���M�4V�F�{�!��0R�%X(i��yP�S�x���P��l����+y�&!||�z��ݜ�����ثc��4r�7/�1���
��������,S����1��S���iZq�U�8�n�ki�}�}jD�q�܅��a�}>��|Դ�=؊OƟF����	_��9w���L]�OkJ_f���#��Z���K����\��z@1��ȓ	�aN��z�՛���c��ї=?�(�Y�5��MW�(��,�Se�{�����w�Tޭ�:G�o����yu,汜��?�@������R5�=<
aF���v_Ish���'7D}^��|���b��no06<�����V��)�z~��TV�t�&l��Y��G̑����q�h�;\9���Q0�;?�(~���tpfw[�tKS�3�eM)���%W`9o��sr��u6���U�֩�S��6@N3)�<lE��kcRz?�3�{x�%^���м;����	�Z��b,�\*�X�X��a��v[��2G0�J�Mg�(:�c�lJTt)\=t]3c���o50Gj��H�ҖZ$ ^�|�9&�f��w$��ܗ!���ꘙ�;>���m�5�ǌqo7A�y'woH	�I���޸�a9���.W�k§� ��6�[f�;vᾗ��g��*��b7�2�h
[d�=BE7D���;{g��*9k�!��J���a}Q�p��� GA�����,�۪q���XӒy��l*�vIU��Y�k����7�ev�V��,�؎n����v��<��� l�����1�*�}�;�ٴ�p�>���oKt��Q0��ܹ�!x��y���O<���5򆐗���i�z|���^k��ϱ�}�$d���^V���%~՗ #�/ʭ_��0V�]� ��ܮ9Un��}�f��,"kRد:�\ ��	�RR,<�聥�V��@�e�z��wt_wc宅�x/`G��܄�_���8t�,F'�R� �ܨUw�������:�3S�:�������%O����
�J�QԒ�g��l�>�l�~�"J����2�i��`�}(^v&���wGE�&S-]R�J��\��[�{k­�Q�����QHK_E�=� �j�H��xj���R�ߑ&Wz\O�;+�/f>%54Lx�a�S7O��T��; Aړ�?xp�%���\ݕX���v��s������w���b�R����w۳�+3�,Pf��Y�o��o�S�xV����0PZ�?L�} ǫnjs6�WZ�ݬ{�(�YnH�%Ő^��{�{�8��@rX��2��M������?��_ٰ����~΀��e/�Y G�}���Oͮ� ۵wHU��c_��s�S�3(>NJgge�?+�{$��y�Zi�J-7�ޛ>P��w^Z3;R����z~�Q�uK����5
�%.
dv���q�����P-�k���̀m�>���.R�ީ�W�N�~yA���B�iќ�����&G����\�ע.O-���ks?t��5xj�2�j��@�NN7מ�¢�#d�ʻ����ubʇ����.՛�����O �<�G�����.
a�#8:��;��bO���ы�m��kϭ��
�x���7����t�
n�'nq2��S΋�j����ğ�����l�b�t���aR]�Q��	k��xϣ����s/�������?��iht��4(.FFx��a�&A]h��uG��5��6|�1b������s����S�9�|c���K؋��Ni�W���94���"�-Q���O�����P�NO�;���y���kf���E϶���v����ˍ��ޱ��U1v��ͯ���d�]�Su�w�#E����%�S2ö=�,ąo�1�4��������<%u������Eit{)�VbE�L��� ~.6��L��y�aSx|�����]���x��|�~O�L'vn��S��ׁX�H�k�������P�����X���U���8�;T���'��[�Y�q�4��� �|�YF�������_�n�!� z�ИQ����.�Jjũ����֫P�����Ώ'n���8ύ�o���7�.v*l�B�Q�c��[�+�t�}�v�x����ޔ=)l�j��`��i�`�u��PY�`�fd�Wu��s�=��l\ǚ�h�\I�up^�s�"2zY����FY���ˡ�������|ʹo����A�3d��o}�$���^��ZVJ�;Y���PȪ;��.sG^E�pG�[D@���	��ӷ5vZ{i���o����||yd!�m.S~�B���b�C56�>�g)�7�߽��b5R��>��\Jz�%P��]}?��s�jbK�F����>�4^6�D�m_�L�ۋ�<�ЇiZ^h�d���v�>��9i��͒�no7 ����9�R�n���&xҝB���}~��ܯ����&�e N��mQ�����&*F��Ⱥ��m�O�s�%fI�}�ڈ�&�ḯ7(�}2u�@-W<3+�x�5r#�P�Ԃ�i�!�\C�gC�'S�J��Cqt"���f���:�b�U�ӻ�E�B>(�Ӵsy9���<�V���;[u��m K�����=�0�K��>�1�_�2�=.M8Z�\�Q��!b�T� �ki���S�]�H�4�:�7"��z����|���U$�QW�v-�I�� ҽh��g ���S��u�&�gc�l�Ȥ���J4dE��vcPܝ�dpӖ�"�iM�Pa��6
��f��ATB�����3��OFj<�റ�n�&T���0�ۺ�- c�fN���>���R�k�jXZ��T-��l�~��m�!��]�xH�o:�	����.�P�./�t���lњ��ZfԳ��&'<�:��p��Y9���d�h-��u�E?�Ʃ��������o��N���i�0��/آ:���Y\g,���P��%�w�f���n�c"�6����q�A�i��������Sn���!�TT�,2���d�W�e�ʲ�'����
B�P^��x��;��������w��"�T��b(�ZͮNR���ǖS��V�nT!��i�Yʕ:��>��DN�~����z��ј��E����a 8bl�Y��~-[kӿ��1�
(D�d�<�]��2��P��>=`8�'�N����"�̬��M?��u�>{χ.-`R���jk�cA��M����i�e�Tݷ�&��o�m�]�r�	G=�.�����<�Q�ͥ�*{�`8���ȈY��g�rոA�T�c��[�o�'{��h���o�M�>�xw/�Mꡑ4��3���8�ڠSP�ׄ�1Λ�L&�/j���jx��&ӓ0A��~��B��s����X�\��Uޣ<����B��z�f+E�j�oʹ�yw݀oy'\�8=|����,�9^��vJ����s���pf����8�d��ח�-SIb©�����$��2!�7ho�L�ɡ� �+��`��Ԛ��'�L��M�[(�}���VD����E������q��S��ν�8�	7^3sd���4Ě�'ЈmD5��>`{�҇z	(������e�!ʮ�ľ���l���``�"����[�} �k#?xpayR�e}Xk>�ܟd�"iD_9�7#6�g�.��}[LVy�ɢ�a�.o�m+a��xl�f@[vmz����NM=vD�#dcFǤLJ���ʦK�o���iut��Yx�Ǫ��4ҹ;����0��."����K"�{aDU�75�ث������PiL&�h��	�6��v�`��'_
��\蝎����bє�^����U@���^�V|���Q�u�yJp���M_�[�c�D��
�[�˓q�c+n{Qx�t%t[h�=���q*�p^�]1&���%vP\3��@Ĥ�Y��U8=�Ң� �g,���ɉ\�������ݤ[��QG��v&�o=�=q}�Qs�޻
D*~5�M���*�b��u�u\�~z��qBt@� �f�=��ׇɗӒ!��jZ׮|�1��m�z���8�c��Cz��9 RE�������#���*pw��>}�±��z���������'�i��}��_o����<K�dP�?˽���9c<n���?�|47:��F�"㒪�%e'⧕k�kY�&�%|���}5�w㿶�o����'���g;�sx�t�E]�H��9�5''��}�a3��U;�N�@+��#{3�:k��?�4әJd,�����	6�5_ �4J�1��K�j�9�*����zͫ��t��Z	�m�_#%�>�T�{��������H0��*��i��*	���=�U��=�sP��JDW��}�$��l��F���?_+��[���Nf⸮�I�7�n��7���v����`�&b�t�+Յ��Xj�sB���|7������Z�o�0��Z?7�ȧ��4�vDl���u6}E�u˕>���S5Jc��(����{�A�mnH�X;�;�t5�������<J��ӞM�N/V��bNFB27a���:��a�j,E���Ρžu�f��&�}X��]yt��R��8z
V�5��������>������Nli�/�ס�����+J9{�U�	r8��u̞��{�؂_~�b�	_{�� ��:��8�.Db�}��y�NX/kX��f8�-��I��v$�]�!�o%E
�͙����'���4Ͻ<�R�l�jwav�jV��͟����"�{ą�-{x��.N����l*iw}�|��2��dF[��	���2�p]zg`?�zC,�cR8�����>^���L�~�wCza����h�+ι������o�YOjz��.X+n.�&�kpn�IChAR�?MP��(�Z@ZT6N?x��xzBY��s+{6�p��`�6w���[���U�#f8rG��_qF-�52�'�=���ɫ�.����?����{�Mra���NO���;� �6%��uÒikS?^��?h��4�Gh:�On�޲3�o6�[�W'�#���`T?w��/���K�[(��Oa�qt۹���A�or@�}�BDG�σ�@�_K/:h�ݏЃ�[�,J~�al�}��f;��Km7svg��6�ux;�.qu/��'W�SZښZl/��e���!�/�D����].	g�0d?��;�~�����Y��q�(͟�{F��ƀ�����NH@��&Z�ڴ|���Wx�ĈZ�}�1�#b��u�&e	bJ��}k�.��>��6��M
m�k�	��a�w u�s���+�wP/Y�ʭw?gx�����ٿ���$Mʺ��n����R?�`�Y1ϲ}�١�8^~��r���X ��Qb��c�J��3���6C� �K�����B��y�����,��k��wH?e�ʋ��Z��$���"�TO�w-'���U5��ǲg�3觻�x؏K?Tk[w��G�:?�J�������%/l�w����֮������Qp�<؀�d~�:�^��ј��Gm,U԰��
���E�������� ld�s&\��1@��6��e/���^y����k';�,�S�X�����iS�������_��>���X�G��h���PX ������ƨ��p�6Փ%'����O�B*��n1�@�l�����O�Փ*��`��	��,���J�^�/��L�R��h���ޏ���H��Z/w˷�Y:�@n�
�a"$�{�Y�D����	�}z��QBz�P�rC���|�mqB�l��^�@q��o�8_hF�x�B�8�LW�FU�im�>��L�q�[�%u����@X�	��k�x��Ƅ�5�EæI6��Va՘��-h�X2]M��Ѧ�a ��db�_��ŜMh��a��0]�wGQ"S7W����
��_(�|�hOu�NS۶���}�F�������`��K��g�Bkl�!wsX�������Hu��h�!�6������!v������ӳ�oaR�N�ub��IQ6��,�R�L�ε�=�����t[�S���c��_{�!��$��M����t{��=�`zw�Q�3��izR) Yu��᳐�!w�IT>��np>�P�3�s�Js�XjW�_>;0*e�f-޽*��6�a8��|�*'���y-����W���HE�����م� ��5�%Ĕ��h���LM���b�YXݷX��d柔WQn5!"���i�ܽ���kZ��n�
����k��Tlx�p��#~@�k��p��R��{�Sgg�i㯏�]":������˲]�bМ�����K��c����`�l�=)�t��i�\Հ�^y'^�ŤT���qnˮ ��L(�B+�pf��������Ad�O�85��C�:'�p�d�R���P�������Q��Ek�}ȫ!SI�\2[�-���.ʋ���!������ԕ�W�z�����'cj�_�ׇ�1^2�[%]���Z�/��b^�Rk��W,�=�߃����7�{n�������~������)/�|���LT�1;A{O�:���"�K}�Pʜ��K'���D\k��'@ؿ���sl<�O^",����7q������['�a���p�+L;���Gp룙�)�d���^�s�����%���ib���A�*oѯ�Lo~���4�k�	��U���8?��W�X(��=��Ş���!����=m�b��׾�Ř/� y�Ͳ{��ز��.=��^ba�K=�m���!����]��t,�ӎ�W���KzG}�.�he*nۂ��F��l,Ny�s�s���Oy���g�?�Ǐ>�����${3�@���Ӡ����u}:� �'�u�4���X���o2�<<jS�ZS�v	�x)�W_~e��mo�Ʃ�,?}����y�Efu�SG/�_�\�x-�k<�(r�W>b����_rҭO����*�s��Bq�չ��)M��L���l!�_��(���p��|ׯŞ�s�o^*���[��]�J\z!���"�\���I�
tlc�sKoݺ5:w[�S�~t����n����bd�k�3q��S�7�q>�w���~��������[������帘��˯�8��#�?�|���_�����ws��o��of	ջ�;���>��t{]AG����Ȅ�$���8��G?:�����s��zB�.d�Ui9P�����g��_���?��᷿}�ȋ ����c��A���V��5�'O�OႹs�B#t�s�u<��UP��� d[/l�\�o��z�R�N�g���tB��,J��Ry<�p��G}���r�̣S���*-3�jB����y�|��r�G��g�p��ˬ�Z�nI��蛳N�����G|�LTJ�E�G���\p����tW�|������ʮ����9uts�0�~�p�3���i��� =Lg��a���|���(��H�<�Tdd��r����g�^G��,�r�+".�D|Ï�#�ҥL�t��u��(��fl���l#Tݙ�N	c��l��ډcu�x򅗹�=��ߛH�(�2�r���w@]�b�OG|UM��AC7 |s���t�P���|�ǅ��x�sW�k,�������_��.���ε��R��U':Wy�=?ƛ�!���2z_LÉ�S���r2�֥��˟�<��w�n>�������b���˹i���q��z&ms�eS�3�m���.�'[��x�P�z�����{��>��5��Oi16yrǋ�����ƪ��*F���d�}���0}՜�$Z�/9g'G��2.O����8=�5߹��N{v}�7�I��n���~�d�q6�X;��>i�m���78(_r�e�{H7��>n^cy��&��#�n7͞0t���3y`S&Aj>|�=�F�<��+l��y��ĕ��vL����s-�5��k�M2���(w��:����W�x���본���B�f�����}R⼁pz�G}�7�~�=��{MR��j�<8��z󭱑L7._��xӎjA;�'����]�������,�g�k��c�Qlz|�4A���sMp�������x��X���;�t�I;�'.� ��eQy�+��#�����K3���1�����#]I����>><������^:���ˇsW2�����d_'�&�f�1�ý=&�ʭ�������~�V�f'�;w�θ��_ɍ�����������_>���|G#�{R*y�:���Ѥi|�z�I̽��^�7D~���¯~��~-��=���36��ާ����~�T���?<�����3�������H4���PJH��q}�{ߞN�Nf�����ߖ��!�����x*̪�ÿwP�*h�π;x��.g@�`r3��7q.�<��`�W^��9]�[��/��GL�'q��$�����%k�tUN��у,�]�U��X�8�:�
���[���5:,X����{�����bOG��Bo��0c{����;��Ϻ��_���h�<���|�G�{�gxG�0�_�:��苵�Rf����;����\����n����d�.�tZ&qbù|A��#�kp�8��w��5��.�U~��23_���Z5t-������1O(f7�uaV�@���>�u@B�s>u�-S����Λ�9yS�b���{��OYS6��:+����� ��|��Ӆ�˯|���&T��Z��P�Ñ/X�4��m�\���Opgr��gt��i��E��+_r�m�р5�<t��J���S��ď������!�u|�0K���6�`�ϒ�xxxw��ڌI��&��<�md�67X�����|�Q7�bYݹԳN|��}e��u��c�6�+\,��|n���J{����w�Ozɝ��n ��A�?��w���Ph#.��H��p�!�v�v5F���H������ ����7/143Q��<�<o�����������$\�v\�v���^��������7�{af0�������q��H��&^:=����s��2m^Y�'�n��c�a������x����S^鴃�����<|�c>���{�wۯq��O<oq_8t�{�)�6��p���K��dk��w^k�c�tUZ�$έȹyn���y����6��wb�Q�q�$�WV�/��$k�H��-�t�I�oe������(�`HF)曇")Mr)���?rCܛY�TN0���y(�����)$��)o�q`��i��Ҋ����y�ݸÛ^�p�;�����p�:�N�Ox;y5:���<�O��(��oq�i\�.�W
+�_�cB:��6�"���oe�ު�~���Sn~�+��_O���xt]�r���_<a%���58���M��*g[N=ڜ�����ٳJ�q:��
yy���oN�O��ʕ\�w�Ҵ�=#gO��1�'��ssڑM�g�[�jb<��U��&�� �>_��Y@p�5s�p�Gxc����߽.�o�EhSP��jYc����N��?=x����_�a�ƓJ�x���@)&�c�O�t	6�z�q�A:���_�pf�sq�t �X���(."r�Jy��}���b`��Ul�M�{�e0ԆāO�2Oю§s����8���C0a����`C��uQ��@��ћ+W�-r�_�Z�c�a��&1����X�/ŧ\>��SoUǞ�����ӭ��Q<(��X**N��`l�4�4�nQL�0�s���ɨ���F�
PpԽs��O��l}G��kS �<�4EwJ2һ^d]ʴ!t�t���S��`0�:&rT�(ѾS�l����Ӝn�GH�&.儛�j���e�m�s��lh�@��� hP�������w٨Ək!(N���/��[�yx�����<N����
���~�`l���#?�����U��S^��c���]W��#(�v�:��:����fw�`4��ݢ�;�{�ʒ�j�h�o��N7J��(�De���
4>1�#og��ڼR�x&�X�
I��G�����LT Py'j(Yt�t��>�<([��^�H|�x3B~5
K�g&�rp
��}'�Ȇ��^�\��e�
���y�S3�VQ�ݓFX�=���v�V�)��]8'�Iv��w���Q��{E�l�6�&��	����pw����6H�H�Y���UV��A���S�h�W+iwh��Y�ٷtk<|���
��K�o+>��y�CK�������{f��'��.���oD���=�w+� ��F۵28d����(�|+���9���¹��=���[ل�_p�7���m�ޚc]��uusk���P�g<���pC6c����j��DpKu��e(g.�[X�{��H9ʩ�)�.S��{�5w�vˑ����U�'y�UM�������?X�iy�-��wM^��I/��X��k�/�X+�����zE~ߤ�I/< ��u1;ٲs�A�$/�=&D�P�Q̀'M�W�
�<�n�Lj����(J�.h���~1�#�o�bsN��-��ǊW�Z,�8�܄��}�|��<R�)����8�Dz~U�Y��!��#����j�Lv�7��@�I���G}R�(�&��8��zV���a�o:����lh��w��Q�uk(�`�������8��������I:4��Џpе�?qgq˴z3K9�iqK6e/g�������uiG�kuhl�>0��S�-��ַ�vh�Q�vp��(c�=л�o��r[��{���t.�}����K��%�|K&̯mπ���iמ����G9>IL>W#;nEV-G'\>{czc���wޏ��Kz���S��gu\��(YrA��c�f����S~<мQ&���Z�螪���}"wi��M�K�O��@���w��S�vo���T�S����_��z�}��F�F#jW����;��)=�`r`)�;w!#�S-��iђ�gV@���
��K8�ٳ[�pMX��5L�Ay��fH0��]�N/��8q�"i)mVkT��WrٟtҸ��������<M���}��^%����t�҂9��Y��s��b4|��wreW?t�<RfYV��ذ�\�l��
�#Y��c*y#����J��R��D)+) ѯ��(3i�:!���@JYı�T#^�S��	SG�<�h�t�=9�y붱S��ʡ��Si=�J`�0y�S���N;��w�TT��Oy8~pS'lE�G*�,����j7xM8Zy+�<��o?�ߞh{���V��:JH
��f�׮����Q�����o\V:������Z�ٸ���#0(]`�9ah�ܵ�K�}G'$q�1ѳ'�7?8s�9������}�f�_|��8��N�Z��f����N�PFG=�V�zxU��m ��'���mP��:�9&��5xX#[�[!�x���g��]]~�M�(K���-@��RB"/�x�><�\�3c?�7l��3���tjل����`�B��j:����;8��O��בǠ_��7��uM���i���ߎ-^���+9A��>���W��y{��y���l6��
��w��S�z"�*��	����ߕ�,���o��RAm�m BA����1C-�G��`5q��}
��Q����i(��E��[8���Oy�q�ȇ?'�Ap����n�m�̫I|&x�k3|8�LX�J��o%�ˉ�70	<�G��#wĳ�T�tqp_� �� ���6	ߍ�t����4`��o�i���4�-���A��IY�<F��K�T^�ȫzL����2�@79{�l�m�n_v���J��<]?V������4M_<m�����0~�Om�?^ݼeO�9,7�M���X��[^�z��}��pտpqq���m���s�.z���]8�DO�-����i㞮_��9:vKNNښv�~��t'3�u�o�\8�e���I/�o���Wx��[����/39�8�i]�Z9fYN�#KӚ�o*������Ӷ��G����*���2����=1���ܖrn�y:<�/]�n�@����iu%'LB݌��uo�`���=�*���2�=�7�>��_N�<p���>�HY��u�篇�Ќfid���7b9>���~��؃��V1�ފ��1��/�Dpi�>�h�̙3�8��,�b�ZOEo�+f=�E���a��X�g�x8���l*o�����`��CY	N��fH�O�@8�r(E~󟯸N��p���������̨pے�ؔ�F7ȅs�U���$7F�um��,;ʍz*�H�����F�-�QΠ�6ۜ�T'Q.@�@#{?�D�,�"��D��$��ꄣ�օf|˗gi|udfu=�z��'��kY�j�Nk�.�E�R����&�ss�6���Su+u (W�9��Uy$o���e�)(	/z&�]:6�-W++>f�ƃh4����Dt
�F��K��Dy�˃��8�2�G�W�<�_��)�t��=f�m�,����Ԕ~���:�+W����yÍߵC���;%�����n��������Ɔ�SY�QO�&�[wN�ʛ�N�{�%�Q�A����+څ����0�_��/N�	̆�
���ũe��"(r�l4�['U
��(�^>]�������p⽤�2':�д�%�LB�n�nS�j�o�JQ\����
����oNʔr�Kf65�����Q>u���>n��Qe&�����^>Mۊ�?��M9j�3�f M�Yy��QL�D+�؃�iG���1C��&��oq�(���B��
mh��u�ܭ�2�_����]�R���V����]�C��������1�}�S���Rx��ɁQ<�2̢?�kZ���5|8��0�c�.���VO����N3E�R
�/i�d����:����-��p!����7<6D����!�8�m�)x�Xq��@n>�_�i��&e��8��bF
dn����`���l���
���
%��@~c��i^�a���_�r{���g�І�AP��\�ʃO�D��Ȁ�YT��n������k++K��q��������N�]��&c|6G�����mg< �^M�,�3�t��Z��F�'p�&I'^�%?0���s3��P����twUl6	�9�s#���L����ݳyڔ>�����`�V�������U�)�>���a��8U��[�r�}�3�ҷth������Vr8έ���ؼn:�pL�"��ә��|X�qn۶.��e��c�b)�����	3��;�P2!ta�:_���5�n�y�W���u}��V�8th�n�j��{�(��������ȿ�_Z�P)�N�jT_�җ����/�(Yc
�
�{�����o��1�ՠ%�;��1�8w��t���������0w!8������
�٥A@�(L|;di4 a�j�04R��K;��M+�J:��O^���f�}	Ƀ?�*�o&MV#(���?�PR�9�Wr�t�����sc:��W0��ì�@%�pf=z�c�zx�R&��ie�./0��Ol�"D�ǹ^�>��M���R�4��e���mV{��,��G�h�~�'bqx���à%�a£�Ш�t\^����'4��?\��g�ý�%?u�J\��Z���ڬܿ�[�����L~렸���͒x��5��m��5\y�������vu��Ŭf!�D�cR���GQ�(�L7ne���8h�������.M�����<=�w[�������:~�U�O�~���H�[��I��uT`�thr3
'\7n�
`5�*�&�:ƪ�]��)
%�YshPx�����(G��W�C\���F�d����Ȕ����+1e�4R�6�<ڐtɶxL9�e����jg&�W$-{������uA��(8�������N|aN��M��߅Oh�L��*x�Q�)�g'�L����ơ�z�f�֡��+��`v�	������Lp�Q�m�<~�'e$��Ó�-�N�x������������{��Z�e\�%^;�`㏥\v�L.�Dw0�q'r��{k5�F�H�ɿ�&:����۷�	I�^���G?G�����\��q��R��-]�7�Ɖ�T�!�w�����(��ڧt̜�U{�[{Y��@%~�x��CO���Y\� �oq�C���X��0+�Y����dQ�$mE�~����+\��0~Ms��'��+�n獣8��<�����̀li�<7Ǥ�!+:�[{�o���ԣ�S���V�wN���;�<����8��%<�E��3�_�n����8yw9�j
'0����f`=$�G����Ob�����DE,O>8���s���9m:m/}A��
'
�� "t��dV��
�_����m�2|���6m �?�(���¹���/<3=�өv���T��8���ѯ�F+�'$��n���G2��B]���z����/�G>��W|OUB
0:��W�Mo��nu������3�����_�t��(s�j���a�r�8�Dq@8m7 |-m��9�K�_��ܺ6:Qp��X^y�>�;�`���[�JCI��H�����3E���E�B�G���LW�7��N�F���]Z8���L�Y�2 �-�*c�O�2j���E#,�^�J�F��S�]�\��@��BA���5Ӥ�+Q��/?�Q�(po9~�(�ߖ�/]�X^Yz��i�4�+�f�w?�:�7�������(wZ��8���M���o�c;'�|�xJ�t�:a�q�����M�W����Gq|���|�i���30�GI繝�0��M陽��cc4���x�������}P�������+m�%8~�)�ߍ�7񸕘���z��F[�k�&�wz�<�Ój0�c��k��h�8�w�:�1�=p��v��ԝ��{Ĺ�`:�HYj@Y�&x�`����Y;Y�T]o%��ȹҎ�9�U5h������w��������Gvi�~k;��Y+��!����n~� ����%8��op���q�Ev�p�lx0}�����I��x�oR�2�<���ה��{�Fq��|H�(��nY�/��WzN:�5g����c+��d���h'���x���F�f�_���t&Y�Lҡ{;��ҷ뼔_\fmVJ���p�Ǜ�
�^.�`�p5&��S�Ī=-���t\��opk�+���I?���Ql��@��I�2�0�Up�7��/�ˌ��:n�O�A�hQp��PU��uI�7K�y�0�R�4��=C�=̊G� w���{�ow��m��eh��Q�w>}�ǘ�i3�M��I�[�~�o�M��[^������Im�U����o�QOLs<�M2Hw}J�4&���7�-S���;�{��#{V3��.+[6e�ř�Ө���?ӿ;Y��'��9y�@���=1]��7Y˷��H��`��/����ӎ�I�2A��9���t��2sZ^^�.d�ǔ���3|;��z��5����6���pB��[i��γ�_0������A���5�+l���9�����瞊~��!��G��W����w��J�,�k�r������6d�ǹ��x��7�����������*��W��'|R̻gϞ0�8��bVNzp������G��҈|���-9'y��\a�B|�! *,yY��aϗ[��7��f�_k%^�Zh�/���޹�9x�!tK��U�������7W������l���9�x��q�q���q�\�����v�׃w(:~:mx�������"p1�|/�-���ҴpD��B�?	����z�q\n6�m͒6�i��ߞ:M!��S׉�v�~��O��\���������Yu���S���VZ����y|ŧ���mp!/�u4X�Ɉ?:K��?��x׮(Q�%f�NXQ�]F3�k.�
�ٛ?�3���<� oxd�ۊ�ۦ�!���.������h-���o��T^�������a��[�'�`���R�,�*l��'�V����ު�MG����N�u��sҭ�;Z�p�|�#oT�w;�S����׫[��q�|8��p�2&ͦX!���N�Y�@�f2��m�C��z0��ɿ嘷�5��p�w`�	.>|����t@#��'ߣc)c�{C�S�p1ʣp� "�^�n��o�G���z���A��k��1A�L�R����*�vT���:����:��A�3�,d���K׎��6�?�A߻��!��ݛ�ǣʐ0oeD;� ]����e����w���=t��d�IS�39D��Sv��ZW֍�O���s�����U%�o��-�x�hX;�'��crk���<F=v`D�T>�j�mv$�V�KFHϤ�c$}�m�X���q�~ԓr2A�r�R�c��N���u��S�~���m��[�ɩ���y��f���:�2��YQ�C��k׵�����a���cF˔Y��0�k�"W|wY��t3�~�	�G+V�5��w쓉|�B���4��C�y��ty�ڴ.+����zi%����;M�驊?��<��~�u���2uy�����oq�z'3�̸]%����ūәs����>�ۧk)�M{��,fŁ.���;�V
[dO?0�Fd���4i��U;�寬���<Ѫ�h���B�31u�W����v5C��F��KW@�n��픢��I�������z��`��X�;����W}ϧ�o��üI����j���0�<�U����'��`"�tJ�Q�������!�o�>q�Q�ɻ;k����[�~��n�yH�4n�k��I<����{�7{��(,���݄�x{ˣ�O?~���q�{f��,m�`a%�IN^pz8+��ț���ȕ�4���30RF�i��LϠ۵��^	�8O^�5��#I��(�fl��do`˘YÅDVB	��[�m�xW�ܷ{�t��#e�~�'e#TK9�@�����7�W�2t|����=�[�s��N��'C�
�u�ԍy��'E �9�ҙ�L϶D!�x���W��<.xc��q����Ax������� ��l��v������(~/主̺��,I�D����2�m��YNӛ_�\��{}��[����p߷cj�.��O�K�Ǜ?����S�%��VX+��7.��O;�I�#Gb[y�X��9��.S'��v�ꁃ'��>����A�!_6&�.G�� ���l	~\�uV^a~�P}T�x��u���郧|��̩�5�
�bv<µ�N� �=���|1�YZȠ:��lrF��.3�n�Ӭ.��en�#��9R4x�7���+�����z����[o�}�������u�g��V ��WG���8�s�y��h��I=���sE�?���L�ӵ�x� G��"��i�4�Z�GǍZ�K��Ɓ���&�_�l�o�:��`U�o����j�rC�n;��l{4�&���9�Z�n.E�x*�'���B�P�Ʉ�C�?u�{ғx`L�����ɯ_��wbT?BY���_�1y׵:J����?#�d��a����P,�Ң�W����
�����K�w�o2_~ҕ�y���$�o'���V�E���9w��o������]Y�#�L���|��x�|�W;���� �}�ǥy���0�Цu����8^�<�'�v�G���N���	�M1���yu1�I� �s?k�M���`�-ӱ�7��7�);S�2�\�� 4P_xZU���2F�/�ų�l~��]7�u9�A�A�����V\<k���M77�n��/E�x3�������+7"1di���@2�Mm��lږӓ҂�Jx5�
�8�&��s����r�C����G?���̳OMG�<\���u��.[}4�~��'��q ���A)/�N�����*����_]k���U�̫�
O�j��A3�@��w�����צ����(ۗ���[���f��E�p����Ɛ�����ء+<
e�V�tp�G�����w��̬x#}jVI~[���r�&w��8|X�\�7�>p�|��c�%�t�$�v�Eu
I��W6G9�M{�c�
���@ط*��YNp"ak�\l{��R6�lH�X���� ���Fzʏ�����덜�e,���U��f��Z0����d���'NEX�.!e@�np*��^�FonͿ~��W��q?*����Ng��-m�͚ԗ�������!]�"p)�h�A��KY=�����K����[m��v���W^�^���ɒ�ѣG���?�_T��lp�ם�N ��q����å^����4�
���R���v97keb�囥���l~��ߝ�}�����ʱr4}�\�18��7�@�Y��g��󆢊����ˊ}�~�`�������R"����կ|}�o����^+���_�z�|Z�X`p7f��푏��78�������Ez*{"���\
Y��t����S���뉕-1�ٻwugϾ:���5٣(-߼R�V���{ ܥ�[+
<dՃ�T����w��\o��D}Ñ#G�^?��K!q�9^=v�X(Jh
��>1�ع}���t�{�R��	�Rd2c�Q��Px�#/���8����o��hO��������k�-(C���.]�Zm�J�4�0D�4-"�����X��脸~�_J��p�i�����enYв���.�"<hA�pڜ�j�&�#\�f�ԍ�g�;.�<�%2\ܠ�F'��IE!�3ٛ_ɦp�r��J���<��$˘/�I�҈Oqk�f��2���7gF>����l�jT���3\�&�l@9�p��%���g�O@\�_�u^]^�vh:»}�ރe��+��ރF2��9x�`&��Ռ�-z��8�-/��t��ɳ��~��p�2�#͍�J��P�ՠٸ��@/5?7L����a��>Te��`0&�1�M�EDN�L�X�u�r���[��B&-���0����4��溼��?_W������͉�t�]WR��L��C۰����7^��~Ã앻�Д����r���h��U/����;c�-7t�6�&+z����9��LΡi�`���'����F�	�2q��>aLOL�_���Q��T�(�,�kT�K$��9e��g�2��t���<=F��**��v��|^�?O�J�M`J3v�����.�t�ҹz�{w0��y4�5�t�~��0�ޥ����|�e�9����S/>�u��ql��p�ظƍB]f,_l���4P�x�(��|��Q˅~5$��	�d��iA�X���s=�хb��|�0�e&F:.�b�����[wg{���92�s��̲I;�CfSu��,X�J��Y�f��Μ�pp��5�W�D/8,����ً�ȓ�ǧ�{������=|�]�������a�߿;\��[�jP����o����?��?����#5{bS��t�R�Rt<y�����o�2�WZ��L�V׷��(�Q.e�����7��'nߜ��t�÷�cF늫	�6��Gy�3K��OD@ߘ~��O���?U^`
�W���c%l�.���1�e������ ��LѲ*w��C�v(e�?4��	v��~�ӗ���?~�+�����c ;=9��XL�b��hV0rX�ko�5������M~\�d�=�g�l��G���oB۷2*�PufCi�ǁ���We?Ԩ6���攞/|��cO<^������{mN�(_'Wq6�_��4(�&2�
Y�[z�5��3f4�ȁH�J�Oӹ�	����QԘά���~��镟�<m���]��x�rn���}��{�sqص�Ӆ3ǧo}�;Q`�d ��,2m���[��Yf�sZC�]��,��ͳ��z��*4����L.�]�0��k`�օ��(:&Q��L��}`Z̪ݫ��\�>�,x�x��r�k5�A�N�I_�K~��&y�*�L�H���M����]��ׇ_�$����G�>:�>s�xfg`��ҥ��=���O?��/2ȺU��~ +�7��c?k�	%����V�x����u���u��L|w>-J��LV����mo��
�����"[�A���-+p�#�I� ��dS��'8�c�Aʄ��_�C�҂�M�/o��+�>�5���`,�+xC��`,���/>x�NHw��`�f Z��:=���L�E]�,:�h¹�o�D�4���v������w)�j�gn��z���yq��:�1�ʀb�#I7o��B[����n�4L17��VnG��3T~��: ¦b��3����U�
����XI0X�l)^�p��t�����+�k@?����R�WRW�c1Vw���2�����7s��r�٘�m�G���L8��7������-+�a����6t����d��pK=׹��D�:I�յ�����.�;�iu��k�4�K�����]a�?��0w]��[unR,\2]N��cR��i.�Ϳ�;���4im����?:l8<��9�-8ek�����נ{)9'�J�e��m���==}������	x�N	�I3��Z.���*5�-�q[s	��O?]�'N�����^�QJJW�Z�t�XfYte�~��Os�F�����|�p~���ͯw�gL��:��i;�ǽӯ}�S����u�Z	�&�u��(B��_��ƄҠG�0�0=�lE�_�W��oqN�i|��-��������,c��>ՙ��o�:K�����Ώ��3]?�t.�]P8�zcw㲆Gp�:ܷ8��ǹ������?�}����`k8=`�ߵʓ4!��3���~��'��s�����1�ĉ��;�L��?��G?���-=e�.�Dp�R�jc6�u�-s�l�C�~��o���ȟn�~S�궔������|�x�1{V�?�pű��}{�+���1.��NLx��{}lZ����(���*W¼c�5�f���$jZ�´{��k_�j=��9}�����/O�����5H{��ߛ�����t������c�rb`$O��Z�Y����*��|��V��A)���Z1SD�˥���&���/NO���B[���?��׸�4^�NdU�`���͌����O~x<yw�r�E�����Q.9x���)v�;��s]�
��)m�>���G�G��#G2�|2��D$ʪ#�ϝ?S���jvЊ�����?�i:q��X9���� /�;�A����?4 +(��A|�mz��VV|S��-���WL3�:�ݻ�N��oڛ7T{�g#�����7�9t�^<e�m�~x,�rU�xq&o���Sw�#���8֑�Ν�������{��>x��t྇R�k�_�Q�W�g�}vz晧J�}����w2��^��7R���šh_���'��,:�̠J˰�|��;�!Xݐ1[����M	��`-�W����N|J�MzC`�[��A	-�S� ܓ�(x�:��(G�!+q�����[\2�x;���Wt�9%f��G|+��W`]͌4�q��h�x�~3u~;��fs%eI���fx��2if��ُ�y~��7w��nݵ{�S�sWr��ɝ�wV0�%����n���}G�Rl�V�����dPm�=/�3�P�[�Nv}�_�"�L_�h�� ����g�ӧΧ�瓫�����<O�����b5}��\�|eښ�?�Csm�V&�䅶h����]�z�F�8���]^~»�_\x�����������*��H�q��­�
wm�*��0p��4����t�J�V���9Һ�#�Z�dz'�~��_���\�O�Ѯ˯<M��U���>&� #�3!���3�<S���s��Y��KF���>�F�c����'�?bte��7��[�{�a�1f�9��{b�����0ۧ�.���u�-�m�i��Q��)n���7���ײa~��g��AT�aGuۛ����k�Iq��G�v�t�����=�'����'H�BIX!��p4�%�tN����,o���g���3�~.��'�|�kZZ�O+�"���4?3d�n�(���?����,��}�J���&p��U�IxG��t��t�JL]b�z'3i܂����K�B��%��߽�R�S��gX�욏��0�Cce���[<�yQ=�O�ٶm{�ږ�X��/|)�r������ۘ�|�k_+���?��|���2Eٚ��B��Ւ|���\�x5+�%�T�]pܟz�ʂ���sه�e�������#ܻ{ON��6�^��`��1�����_��K_O��ܷ��6h{w��æ��M�dXA4i�U�Ӳ�YB�h�V�nGI�neM�)��'�A��R$����R���a���]�~���������$
x�/3�x�fF���O�����e�S~���=35�'V�^}���O���Ȋ�b�u���#���?|�xg��;fLk30��|��R�a��!���;�����_�x���Y��� l
��	�-�w����K�)�����Zo�Ĩ������ܤ��g��c�U���n������;�;�� Ԫ���ƄOx���t�Lv��՘���~Hx�π>/Z�^�yW��{��{Q^�eP�՟��Ƞ�gY��V����J�@NjI]�f���ޞ^z��?^�J�oufC�B�-��Ze�Ċs�����A�}Yeb�s�3�}6���Gr�N��ġ���(��2d�_�;  @ IDATڷ�p
&6d���7���7S���������tV�����/�ѮiFɜ���G��k�hȃ�g�ቧ`���\���5pܽt-��q���!5L�\(x��������n�(��X�o��p}.w��}��uGV��N��^��(m��w"�:w�U�q� �Ů��س7�0���={廘�od�`u#�7<s�t� >@���w�d�:�W�:}��br���/^��VdY��}tPA��M�
����W.O�/�L(����&GƠϪ�B����.��>���Py�Q�U�H�!����O]�q'����8o�n�C��'�p�֒��g�$:���)��ѱ��ֽ�o�9�#o�z����~�O�h���>M�\��rEѫ�
����}�ј9=_���?ޥ4���}���	�UDUV�=��׿��꠮\�T�ܒ��1ĪA�!ׄ�J�U���pCZ����p���o�ic~����q�0�o�4:8z��quJ�o��M/�|�1ьM��o�pVw��5��l�+¾ˊ��{&6�~�êr�T��ם�{��'~ Kp��n���G�*opl�ĳ��|�Q�ۯ��o�_���|]�}����{�w���������t`�7S��]@Q3�E�q@�Mė.�,�:�З�ή(:G�-����3A'��N���O���2��N�e��z��	ϧ%^a����N:3�jmC�G�ex�g������#OԀ�	u�R�@=������ߤ�˭ʁ)|tʃ���g47��ی�k��2�Q.~���}�J�a].%Ѐ�G)���� ���r|9�	�J	��i�m����?��<q��CY�(;�>�bC�RV�)�O�ط�H�p�,�[�n�|{b��/�<����rE�{��ק�~�B�i��W�T3����	�<>�����~R'D9+]y8�M�kyʗ�pq矮<�ޭ��������;oo��ԩ�Y�9[3��������]�lL�I�o6c����_y����{� +��c'�ס fo�Q(�7Cj@af�&+B#f���,hI��з���zS���~��e�aM�{��kfM���19�2��	0�E��fBFy�^��xah�i��Z��in}l6�����ˇ�N�|�A){�I���s^2��}���X
|��p���[+Eh��f^����kP��F7�S��֬&et��ӥmkR�EX��'�������ˁ�uQJ3�]�U����m|���g�у�M��_"�|�}QM:n��ǀ�_���h�kO�c4�Y<�f����7�� ��:N�5��߶?+E��{��v�����k�F7:Y�^�A��g���Z�ّ��:�@�9��͡���Aԕ�x� ��@��ߑ�Ϟ:Y����r���x���ȩ-y�V���ݓ	�q���/���~��W�����|�葲)_��bL��⮛ѿ��?�Cfj����+ᣓ�ǀ���:L����)�}?��^u�Ȫ���:O�����Ư����ÏS�NK��n�~�����q���sW�o}Í���V7kgs��3x��HIB��o8��[�&��׼��M&���f&a��=��Cu���_���P��.�m��
B�U>$ǈ&[l����\�t!6���2�.CX�����C�+�����������ݕ[��[�t�f�f>�w�����]�ݟ��Ŏ�������h�8�K��:�p��w��avc�������aT~����^�^ˏ�@��w���.���P����U>se��&��� ������Z�	��������n?07OCp:�Σ�?)��wox��w���GJf�1��خw��St`�w�&�Y�F[����g֬���n�l��Ft�L}����)ڧ�gK��գS���C;���R�n�3��<��L�%3B�ՕZb׉��d���x��M�����9J�����~ʹˀ�{t|���<����ޕG�/��E�l�+�\C[���p�_20����s��t��,�3ٱcaږW6�fW���.�G��	FV)��)s�S���:���gVwCl�K��c��M��y�p�c6W}t�gf�}4���Ύ���+?��8_u�,��?Hާ2s�g��?����a�Y�ρ�'��d��N�K�{�?�$q���o�h�?��x[A�d��(��.�6yZqx3��6����Kz��!���-��<�2:n�@�켷=-����ޓ���}iz�*�� $� ��ѣ�腦���t����+���������g6߈r��o�n�
�6mʠ�c�kF�DM�R�Z~Ѡ�W�T�� �*x����3�R�V��;L<�a5
<���t43���=~Z�a?��u�ԉ��l�=��ݱcW)B��H�W��t�:�Y���EC{n����;��_�r���R��n{�����-f�91J��vf�0�R&\4N�=�2�
��3��8�G�b&��y(��l|�	�:f8��[Ty�q�AgVO��a�8i��j����������7�+�n]��',s���1�Vydz䑇_+���r��Jx	�9<�;����W^�|l�_�} )G&�g0���i˓��m��-�\��#G2�iz���2H?����jO<���-�(^���N���Ҵ.�D+$�Sַ�|��-l�ٓ���z�:��ɣv��+�3)Vަ'*�G��Sa���ՙXt���+��];3xߨ��)�tX���x\������������7'���~w:��ϯnUO�K[��Wp����\�W��yH�0Gڑ7:V][��Շ�oFxe�?�����#ug�ª0���a�ѡC�/}��<����7�<���/��a�J9R��4&������Mc����?���c�3g�����ENZD��5��G�0���}>N�l�$�݌�kLr/����K���2tH sM3o��0�A�2���/8F����B�U����UF�#�B���r47���O�~*p��@���#���hi�AZWìd6s�� i;�8�~)|&�����V�N?^�>�O��c����:�O
��4��7���_��ǖ�fL
�eK�)��/3X�Fad���KX&���ڼ�q(Y�7(��=���,P�_{��2a��Qک��M�A�}z��?��i]l���QJ8yP��������|�;�'�>c��띻l_W��Y	��?��d|�[�*eE��!��.�>�S��=�`�ZEa��\� p���e)�)�E�>��35�O��e�L �� �?m������~x^��Q�R��������*���n�F�L��Nf�_|񇵑�Z.c�-�n��q��=5{��s�e`�{:s�T������{b�p!�ZJ��W^=2C�����?��W��3O?E��󇢜?Q��(.+�z�5���޽i/
�2�7xF=����`�{�����z�X1Z�@f`�N���/����2~��T�*�z�M�:x|iu�����������(�����e�����Oӏ~�R������ʦ���gShg��d�#�6��Q�d����?�Ѵ1�m)ʔ2�'�խ=
�h�c�[f�p\�u3���(j�-��jZ�|M�^ɷ"&�v��y��ˬ>e�`�9rdz6Q9����c	�B���Jĭ[7����y٫f�s��M�c�<�]�L�B+���/��bm�F��hZ� +;3ÌGѕ�8x(��)3E})[�?S�C�8� p��;ӝ�urm� �1
s�sT��Ϟ!��L���<�'<�炟S�_�n��~��5�.�7��f8���ʖUW��>r�9����x�7�#��ڽr^7�
�-Ns��yǎʜrW�a�����/ե�wRO`Y�t�������F���\,�<mϦ�}�.��rg�ʝLD��w_Z7�/哞��(�<���{ǧW_{�xr�Ƀ�8-���Ø�e�OL^�j��>����>Շ�P�&�)�����=hKʎ�<D⊋.|Vu6�o�"�|_�1�XīZކ\�(�h�RWq ��홯�2��܆��7�����u��~sҴ~#��ƷÍ�\l�Ig��PG�t���q8V��?�Ewo{&��dVF�V&�b��ؓ�M_�ꗧ�~�K��y$f�[��V���k/Pn����W-�g(($=g2�[�۶o�{����V��
�O��B�rb`�8�ڿ�\~�;�|��t���'�����4�)e'	�m��7q�w�7���N�i�����3,�4��jƳ�
N@7�jH�2˫����="5�3+�W��G�1���)�1�yy���݅7k���������Q�-�oF�5�Ăw?���<7�͸�����op>�5�>)N�������垈�v������[��%~ʭ#cnAYp){0�Z�Sԩ�D���s����9�����#\�Za:L�e�[�3�(�����ܿ?��?�ͧ�ի��A�Z5��)�z�i��'
 ��[wξ��f\�����K��-���£K��ޚ��_��3�W3��t8ۗ�!'�h�6�o�Dޢ��(��k7�.�n(���%���g���V���ޝ�~��i2ӌΏ<�ȴ/
�];�+���VmbJ�ߞ�G���1w�����������.%��Cs+E���}������Iv�9q�(�9i&��U/h���Vh�g���ȑCӃ�DA���[��%��0!ڕ�a6���`_N��Ɍ��lv��֛�������aK�|m�W��A��������˙�je u�����ËhdE�yջ��x��m�4���/�"�`f���� �סRի�d)���H�u��Yge3 �˿��<_�aOS��P�c>KQH����j@
����5h�r�G�^V�%����ܵ�VM�\�Yʹ�"%��)����޷}�t=��w��;�0Н[��R�w2(��^�� ���2�~�0�v:�jpDw��
s��<RɊ��g�+9��ܢu୒��cUª�1����/=;y�龃��w>x}������`��X��Ld���A ��`&�p��5�\�>�H!�
eS�� ?�:�S�\{+fG7����K��E���d[�9���Rє9�r��:w)�ef�u6fo�2����\�ӻ|Xʜɑ�c6hc�������9��]�T�f�9x�ǁ_�2��K��ɂ^��^�N��K^��={�Մ��l�V+zgϾ�տ�1�o:��Ν;���j�q��]%+�$��!M�05czw!�`�ֳ�<31kZI���k�M˩��ԓ��~�&���������ݗ�e`�{Df�o]���ٌ_� ��Ri���Μ�u3o��W�Aߪ�C;vE�ٓ@^�9�v���Φ��5���}��Er\(Y44qi ���FO �3�|*!]�"q��A_�8q���^r��S�:(�`E?�
��� ��GO�$o2���n����7Zt�w�w�M�5���j	��O��ǳ�z�S�$�oj����Ì����G�.��������y|)#|��t~��G�d��^}�ן���ģ�e@��D��!8y�W��{�K�g(�2d�2���N9L$o3g���W�XŚ���N㻻9��<�]�{����u:i���nH��|�ǅs���ᨌf�Kd ����w������, }U~1�i�'�����u~�G���Ǩ�Q^�*��t�y��a�W�E��c�"�n���o��qC�!@�1o���yw�#��ю���mz�g��g-�|�:��k��3�n��_��]��~ݛ������h���q���-��>���%�ԅ?HA!c����"K)=�����_����o����g��Q֌`���f~D(ʄ����AA� ��).m^B����g?�	R�,�:~x)B�m�������8�(iW�^���\'d#\ZD�e�͎SVZ(�~�~������N��U�~�ܙ(�ϦC|2�Q�ɒsU��ƌ�v[�nF���a�6}BCK�iJ�zr!Ѫ4�z��wrd晚m�|Ͼ��������?(����*0)ؗ��z�ݹM�=~���k_����3OV� ]���K�V:R�2q���ԥA�'�\3ق����&�h�sʞټ���sԥ`�����5V��T���:�����cԯY��'>�ӫԽ�X��N����s;7y�ˣ��w���u��͚����#�r�cȲ�����~�㗊wO�:^
��Ãp����_�b�fmSx��ՓQ,O�/��'�\��err��0Cp�*�3;�9|h �\N�Q?3���M�R�V�G	��+��;�iӱ�ҕ�@��
��w锳W���}�����r�����x+�KFs�/��衟�U!~i�X8�G� �0��~0}�ק?��?��c�ַ�s�^{鵴���e�R.
e)^1��<=z4
�Wku���=��G1�;S��9�g�)cn8�9��t�^�� m�/\�='��͕��̬�޳sړp�1��U��Yr �ݙ���C�Qzk���b�"m��\�w�L/dՈ�	}�c@!�/��շ�퇗8r���� k~Cn%tk�ު�_��_� �tL��&?�w12�!�����`��8ɑ�Tp?�o���V)ܑ�`P�����}�V�?1�6��PT���UW6�_�ѲWë`��cYoZI���Z����j��݌�p`����O=;=��_���>����1sz��b����Ke>��\��W�݊&3:*{ӻ��?� aWx���6����v�L�e�
�z�o]f������U��Y=��~{��󭕓ę�Q<�GWxt�����w�i?q�>�oN�'�g2�JL���΢U��?�g�[=x�L�E���+Oe5���v�}�ρ*�j1����ǹ��|�~\�{�>s@!�G���f�!R ���N����o}�;��攈�p��<ҙ����i8�<��xM�?��G��I�`>����Fkb�`́��k`������5�rP��B�Ug���zRCj 66���!�(�l3yF��C���rqV�4��\{�並W�Ay��Ǥx��a�i�aP���
<g�kA�_�H�Y�G�����	�ݴI}o�5#l>�\��秥��H?s���˟�����D�vi�t�j�I���=J�����&����W^y)�b%+9*v�K9�{s��v잞x�鹧�*E�
��빴ȑ�Ler��Jڡ�D(��җ���7�S9��@�Kp�_gx�J�s�ۙYw���W2H���jj0�ٷsonA�>�>�a����ePs.
�[���̜��������Z)����Wjf�Q�L�����YH��dR�%^kf�w�4�	�Ɣ�vf��"3�O<�D��z=��Ӧ(�fI�'�R�N�=+ۢ�=|���(O>�t~�(1Ϡ�Rl9�m[���k��OWbn��{Ng�A���(Ji�&�Y8tǶ��:�'��\,u��t���t����NGq''�\����k9�3�u[��X�Hc<�X6]�03��jV��=����;�[�U��2K�.'�Q(ץ,95t�
����g�����F�u�X�yD�f�D�\Ĉs�)�zp���������ϧGR��o��f�:t'g�ᅍYi�����6�{��(�35S}#4����C�m6�oϊ�Y�ǟ8Rʶ<�J�\�`,jʔ3�j��1��y3�s��||��W���^��$�ݵc>Xe#�ㅗ�F)f�9��M�߰+'�v���-ۜ\6�%��R����e�8s5{2�ڌ���Ο�H(���J�k'��\&��_�����=���QL�v�!gO��������;����G��Kec۾�s[�䁬I�<3-��լ�lL1oe �i�N}����K��������Kө�'�7V>��8m)6�[�ӟ�������^���,FVm� ь��b�Ax;����Ws�ҍuiù����SY|kz +=0�~L�"z�ԕO�:�U��Վ�g
�>l3 ���6ƪ�'la�9_�Cߕ�/��vz�!+R+��+0�޳:r��t߁]i��[p�b�W�Ǟ~|:x�����iӶ�z侄��Rב�[�nȂ͑3�u�ڝeG�F���Xm,�?r�R�9R6J�����z��Xp�X9S�Z�� �V�A9ݘv�=+&�G~��O��C'1���g���[�l04�q�Y�L���sc�x��C�y|:�U�����?����ڙ*31�O.�'���٫��C�:���<���Җ�k+t��BN��<��qg�������UG)�ۤ���X���?d�B&.Q��@!�/l�o�`d}ǞUG�����(��!��Fő&<pޑBN��>(�]i���{���1�YX�E�ɃU���h�ʄ7�,tgr�l&rL�h�[b��#7|�_��^V�l��2��S��S_�#�7�/�Q`3�C�L(��"�����G��|%kg���}�o�p�e����K��(��kٸ%��Ѭ�=����1q<x���Iô����>���(���lȟPƈ���)��v�fLO�<_����Q.b|��8��(B��Z�ן�))���o��7%���?�C�N��s׶(�G�?��?���o��������̪~�/d�*^f)O/���<�H�g�Q��_�3�qW�K6�JޑY��;ͪ贈�kY�j�}:&0�[��;#i��m\�̂�c���p�
?���b�k�d��_�@)~�Ż\c����p���6g?B� Ϧ��(ۘ�2�0�nOIˢ�9��M)��l�Y?3���ɤ�l�6�w�L���	*V��¢��ݵp4���I��Νo%��nE�j�G�.��	����Z:d��My{C�sU=�q�vl�U�M�����F�ub�SX�]O��xʛ���ك��}a��|���Q�p�7}��w�8�������W�W5㻜+�ao�V��LJJ!	_���ʾ++@ʌ_��;��1��o��𦫙di8q�O�-�۠��wxR��ֺ��v�f��V)��M����⽣�eU*w���`%�H��N�9ӣ�A����Rq����\ʜU��7x�9�6�x���9���t�����C���)�ou�B��I&su�U�L�5�S�7-�L7�vc&!6�OvF�=|�p;o8�^�����i��9��$��r +Tն(o�H�����11�����7�9�;^�e�����7k�|��ɓ���fu�L�2�[z���F�r��Mca���JW���įV�R��	ٰ�;L./O���vdJpOumݖ@��Q�._ͩaY�BCi�wj� e"gk1C�1w
��l�D;��	��u�g�K��O��;���Ye��ݘnm3�fp�a.@�c��0�˗s�ENu�5����#�?s�L�S�Qwf��ѽ̸�)�5�:��3l��Ω�=�J���G�����1ze��;B{�n���uY��4������D�䯕���cv ���L,3kє��%�Bj��X� �e�؋9�M~�S�@U��,b�9V'@��RDf�̧@�_���C1���lV��?��w�a/�b&n�̷�椵���is+��aY�2�;��Wq��q�C�o��Z�!K��{��y��19��6�S�<��/f�f�%�G+�m_���WP����A���#���/�
��ƓP� �8��y�qJ�������{v���^\?&��@�����vD�-e:�RƄD��Q\�x+�����p��=���WK���0�Bf�d6��<�<JaoFV�2���XC��i�H'y#�ٹ&����PT<�i����P�Xx�7�C��Q��o�|L8�m�r�C�X��POgp�*��u��u�GGp�2�7'��O����/�ߔQ^���f^��Mq�g�+���oO�x�����۹�4��ߣ�`Rx8J�[XŁ�:#�)���Y�<����N��hW��17빔���(j6�ڇ@6k��/5���{�M�������W&�%K�g�33�c�m�L]�_NUN]bȸ0+K��CX���s�⥄m�Zݠ�l𙘏\̭���^�Q��_�) ]nta��Fh���[��G!�����d�����y�|�1�i���p�[)�z�
�Y&PKBO񴋅u1݋�Wbg�ń���~�ի��>�*:�	��2������w�h�A����Qv��7^}m������`E���8����8��>�λ�/�����mC���=��	��gr�)Xg1�J��S����W# �S�[=�Z}4O�$��S���� �v�e&W����./3�ِU���f�1%�%�6��k�#?ƞ�l��K�6��ū������ꛟ�@Ι���H��2��j����T�̱����0�ڸ�޲Br%ʾ�"��6~�]�o�kV�	(e6����I@i_��<f����s��L밒(�V-o���]lT��g�vCx4����)af����o�c����Mx]�&	��5�ǲr�!��w���e�s9+~���.i�K5��._����7�-��G�c;���L}lK��jO.�$;�����31���ˏ電�<i/F`5H��8
<�29[��@W�&.��:ж�dAڙA���ӡܯfE�~����dT�H��Sһ�&�J{��H��&V,V�f�
XE����a�r����H�Ͼ@|�Vl6m�5u�ZE��������^�xé�����Hy�э�?������z�/�C��+�C��X�u�~3�iG�����R!]h���T?�ԓ��M�v�Mx/����� �(�H?�B�Y)�����?��M�O��AUy��7��)�+�u�����]�������Y�?��ϢϿ����1�t��ǜ�����X�X��T�/�;�}K�bOM��͙Q�7]����(7�1/E���u�t�7g(jC��C�@�A�C������X�R^�E@�YJJ�+�t�,EF��]oi���-+��?��?��~����ĩ?fڎ��PB��¥�D��$��졓[�������<�~f�t���<f�:��l�A�Z��U���r'�BEFpw[�}6�R|L�HKX{�#O+ �ɺ���H��|� ^�y�g��5�����ި�2������z�������(���Ř]��v�:���%�L6?�ν��\����G�f���[�э	����O_ ��<̘��N��	��o�W2��BO��s�K6��3�h�S�i�N
>����l��7���L�2�������Yy�2g0NIz��q�����K��6M�ς=_w���o��7\��lؙ�W���uz�o�h=t�`ȶl�U��o�����&���o�>��ས��ѿtd��;m+����]8�ӣ���ÍU����ecV��ԴQ��//'�\�I����H��y߱}�̃Ɗ�v?�[c�d�~ 4�x�l�Y�8�m�a��7ߠ��_��TL��h냞�瘜����7-���I��q�@����d��u��r9+*�n�T���=Ӄ���Z������&��!+����7��٘4n�b$���l���N�?=]��W � l)���4a��3�ףH^J]�������ޖ�1�/��c��:�D�Q)މ��;�gh������9X&�p���ﱴG����/�jB�9�]^m��G��3���ؠ��F(e>}Q��)a�䮬8�^�N|0���t��;�x)��uV6�:��M��s)T�E�L��c�F�U��T����<���ĩ����� ���@�'MJ,`�d��Kx�����]_�K��4�w��#�#��ݗ�]�wM>0��߱K�rpG̚����ҫ�1�*�����B�������Ms�N�
��4.�,s�=�O��D�{e���}uh�M�V�e�D7m��u�������( j�
5���Sa�e�UX�$;v��޸]��
N���3�q>)�7����~����Y����nL��7��g�����y8�i,ӲUg���وk��
eJ��s[�R�0BQ�aoq��('��U�:F��fb�����0���(��)x�湄��̏x��.���`(���]<P�V"�oe�Y>�|���,�����~k����?�9�I3�e%|�p�۝����=K�:��(>��rv�{����Mb���tz�͊g� mŻ�AA�-xۄ}&&���@Y� ��(��J���oJ��ʍ6�)/�Tq�3�R��_�9i�^�\u8��2�}�,��`���YR�����ic��`�S�Ί7 _G�M��x�O�/�|�7���9e�L�tpf��?{�b�>�#�4���}9z׌���ǰz6����X������mˑ�x�j%�J�rL�}�<��w�r=� QD����(����Xh�إ�Q���(�ho�8�/:W{K|�--:�J_h�괕��|R�5�?��h��L2>����lm�A�c%{{�:��_��t���������O=�h�z1{}�\Ƀ�<8�y��]�H�E����� �b&!�t}���Ȍ�[�=���_L'c^,f�8��h��ʖ��6����ȉ��^ˠ��a�������1���Z:�\�f���_dO�s�<[r�T���/��Ř�D	u�l�s��1)1h�U�� 9Ҡ�U�t�P ��W0R�)��W��p.�|j��(^͞�D�cj�٪����68޵ۉ��vfU�࿺z_���:��ӹ��ā����\��қo�1��g/gCvN���B]���K+aIV��#��X�s��]��/em{��hS��Ral��Y[<u�l�,%����G�|	=�]���NѴ��h��C6�������B�-��9���~V��%�:��
�J���Ȉ�9��jd��l�w�������b��ZI���3!Vr�����1Y#�I`-S7f�.�sy�]�?_�Zo�O�DC�!��&4���q���۰�������.m����iǾ�T�zß侟�C��$�/��E#�}���������r��peI��a�u�ZY�C�
a �n�O���<m��/���|fQ�ů�x@����7����1�w 'fl�r�Q�чrn�O�8J�:֙@�&�	�!��l߿�t�+����� ���%Xt���3�<U��?���jg��Ǟ�yg�����`�~���
�t� $Ӟ�e��ͷߚ}��>�#J٥�S��� ��$/��Ӽ�ع�[&"дMxi�:1o�%�4|�����К	c��<�o�,;��3g��̞�Yf1�	f=cO@.Ċ]�e���Ө���dS���v������#?�\�y���쀴Lns*�˄�ɕ�Yoit��<�fQ3s?�g�=E��ޛx/���\�/tur�F��g",45�2k�F�pi���ʘVvN�1��F�lμ�f�͘l�G���3������PN�z�樂�!;���{�;=��*�%pf0���O�.Z���R�ɿi)�ou�~���t��3Y?�mCf�T=d��K>xK|G��D�X��۠-�����͠$�#d3�̒��Uy������]Ev�#��	�H`FB0����*�$��R�������)�Ə8��1$�dB腤+��Y��9��+�W*}�>{w��իW��^��W�E|����~_�4~�0�-.0�ߍ�z����1f�����U|O߉hx�S���$�S�tG��۠S�H�������'��t;z������*�t*x�n�������aJ�����=)�ܚ|��f��׋�H��o�w/���������TYe����,�ˇQ22p$����LN�dmzOG͈��-��A�]:g�\.�(Y��FOz�'�ʐ5�d>�OaoR�Z��g0$��2�b���,���ۿ]\���S�?�C:r��V��~����c��R��O<�["*�?���'�]�ס��Js˒$��\�� �m.�p�۷�/~�-~���U��%q:�o�9����.��_^;��#�o��g�~�zҠl�<t$
���/g�|�������o����,K�/�fɏeN:0{���\���Б��=��ĸ��C�2�Yu�$��ϑ�f�6#wf^#�U�|_�� -��k���[�M>�[�4����>2-�Iz�D���ȍ�����Ԭ�N��<���~�����'?�����.��Ծ}�=�XN{���ff,��!���NnB��C�y�g 
�Ò��z&'
_yY��R�5������X���[ٟ����h�#�`�ؕ{L�DV�_Wӹ�|=G_����s���������Ӵ���� n�`�>,���2}O��+���t�'OG"g��9V؀���]'��ʾ�Pi��_Ж�͈���_������q��;�L�D�̖(#=�s��k���J�P*��9c�x5(*���Ǧm�r1d����%��8�������ٸ������Н������G�1��(�G�}��{4�!y���-�[&���2�h�Ъ,\
�����f���H�J�ч?��7R��bNC�ԖI�8P*�RƜ8�WqȒ)�M���i��wީ7E��^� ?��+�ʶJؠ�.�)0�m���%�'�,Q2T�6�YN���<��-��?����K9���)G�J��W��ҝ�Yaཟz�$&�::�ڊÃ��4O��H�t3��%�/�mv�K����B�dFz4t*ui�_8�]7��c�KG)ʲ�G�T�1�G��u�6n~����N\>�(j�P��!�����6^z1
`F.��0o��OP���d�xN�q�Z��Z8֦g'nQ֎��'�o�"ȫ�9�I��L2�I��wU�$n�K8���e&h"��]�ZF�l&��!����߻s��c)�<�	M|��f��#�����=N+1â�7��|��<3K=����ұ��k9�OՐ�g��ٌ�݉R�lb<~�:�@��[dD������z�ѩ�c�m������Y��E)�'���Ǣ ��{I��E��Q�,�����S��K�Y
�p���]�o�$�Z|��p=�9��Q��_�l7هOY�� J�����C���Y�G�?��	��ͯs����X
q<x'1}uլf�wFaϝ��6x�;���RV��Ã��7��&�j��h੥C��a�'���(e.�3#�=X��:5'���W���a�i:b������tp`��UN�!�҆F��&J���6�Z�%7�6�	q��D��X#wي��8�%b���23wpqܾ�GF'5��&�5���i�>��4�xb�ɪ��ґ0��Ĵ�Ν_���_.�6�g\H����FWݛz�=<��^\Ό�'�.T�����2R�]?s�pp�pg�]��^X|��E���.+��B�ҭv��N[������m��f��En�����������r�h��Ƈ'����ף|gu��q���y^{��ŉc/.�H'�`.�<��:,B��@D�z	�+�k�A��k��t%�0�Tw
�_^j����:+vGhބ%;N$��,���J����y^ofP�L�������K����X�{�}��������0�����\�,���lF4�f�/�K�{'lޏ���� �I�,F��%�WN堄� z啗�u4�A�.��p#���v����Ѵ5��y�!�f+��j2�o��#�����Ga��Z�u.���,GC��Vx�����q`^�l�w�ߔ��X�K����#@�����#�֩(-���@>����>�T�	�2���j�4`��xH����"�,ϡT8��Y����@d)QF���d�JW�3���_����5Zl���ʄ��h:��Fi5�h� wc���mz?��e`�ct�Af�~��B��䄲I��fpyղJ�%-�T!�H��G�$�_�$\��7�`�SF���^����C�#�F�]���W_-E��!n�'/�]Q~������\�������'�����i� �fЫ�['��#�ɑ@��?#����Ӫ#������G�|���zS@u�.^̍������.���������+%�*K�t��m��b�̣�R����·pt��.a)�ŧ�K���\��?�l(���E�rn�0��?�QɅ�	�3��{�W��L}3�N��\�#����,�˽:������YK%���ʹ=���;�V�|��`���g����w�W�*�4>�,��ȍ���)��A�z���7��a�rsL�=�d�rF���i8��o���c����S��>��3�V^�|��r���⃓�eXʯF  #IDAT�[�ӭ�N�B��{YZ�|���(���;�?��0|Ό E<�.�ٟ��q3���j��w߮N��B��`J�4޾�z���܏�Yˈ�ճk9m�,�QT4�{m#1�@�AH�d=�D'^Z
)��Odf���M|��sL�L<e����;8�#wS'l�޳�x!3��__��?������(�/eɶ:��v��?,x�gDY�߿�eݗ�ދ/,N�<Uy*m���Y�I�v������"�W$�2?��v��}����Ke"�_��Ld�ɖӽ�}ʦ�,c9t4Kn��ɾ�k�W�ٺx�bջ��>��(��`�ׅ�dOə���m ����U�۪U���g��4�|)��%����墷Z��t����i��͔�{���x�œ�g_<�8�6�~��Π���0��"�V����AN�� �0�}���zN�!�f��R�� �u�#-[���f��í���/F�>�Ɂ�C%�3:�6�#`��y$�۩Sno�,����-�$��k9~���D-��Ҏ�#�E��~�'��G���p�4zK��<ި6�QէO�ʡ,Ƞ��G�ۓt�MK��\���'T�(��6�7�P�'`E�HVyJH�h��9���(4o��OR���6|p�������b!\c�^�	|�Y;3l���ȷ���+����4<'�m���f;
n���v�_��<N>e��ܚ��o���k{x�͛���ˏY���O�v8�]4řiwN���V%2�0��PS�>8����F���
���ͬrm��9`��{v	�v�`�#?K�r�&�S���Oiv��w�����[?.��
'e\��¥ӹ���ύ�O=U)�.es
��Nn�ޝs��=�\�d���>��w#��v:%�.N�z�f������5�.�|�3g�G�`wηY�%-�Ⱥ�͜�ay��K��xČ�F�D�b��+W?�xwF��郏r;kξ����ŕk���T��4�9�4�]\��1\eƄ<��W��'�I��.L0ʔ�C�����4��on�g��,�Ou�J��.q1��,}1d����7�|#0��8�c���ӧk]󍌰���@F�-�ؗ�zϓ��>�4g�������?�Af_��Q&qR���SF�/~�q:x��Ȭ��BJ�Frw��f����!ݬ"�)����e]C�K�tƮ��{_��J�O���9Bu��ō������,�k�u����1ۢ�ղK񑟸�ܔZ��>���V8{>K���\�<:��������|N��hh7zkv?ne�I��(J96�c����5&/�M��ow%nGq�P3:i�d��_���:y���{�Q����'��}u�if7�A��j����nJ����d��B�s5y�߅m���&�F��:X��nf��^8[኏�����$k�?X��g��:)q�������x%�������.��M؟�������)`��?������(y��`fʞ�H)Qh��Lni߯����dbOxu3�]�Ϭ�痯.��'S/�ߦT*y�n_���eNe����^<�;=�l��7R�/�lƽ&��ɓ/��K��܋c��na��ߛ�;����{�7��_�v5#ϯ�zj���h�̩�(��ʌ�$���w�!�D��y$�S����<�yV�W^�)u���_���W/�,�v<sRӁ�@:U�r.��F���(�O��L^ڀ[{r�Lfn,w�q3�ڡ�(��/����t>Ï2�]wZL�Q��H:��ݦy��j����~���:O��,�<�C鰞O�����\�$�::��T��uz<%CQ������r�-����ݢs��Z�2����J�{گ���ǻx�������,=�=:�H+��Q���ǅ��}O/^z~����r2Z����)z��A�Ң�߉'�L7F��� ��,��L�l�3�䒩8����%���`�������?�`L�BD`0K�:�j���˿T�RCq��G5�@�J���T��:��;�f�s{�le����������W�e���w��4����Ł�|�_�����ݦ���ݽ��������|��u~%l�W��>�GM�����tx�)�S����[��~_�����w����0��,�Ӑm;����~��ok��ݛGEj�ߚ����;:ڿ��qݽ�DIq��QE�Ϻ~��[o�U�	-�^XFᤵ���BUΜ�c3,�9��HN��ӻ�rٚ��ۈ��)w��Rz�7�R؞�zN�t.����g):?T���sck�Y�Gr��R�T��}�n��
\�T�ST��g���,�aZl�w^�]�w0#����hj5bn~6wJ��^~�T�F\���6�)
x�'�{�����F��Ց;{6�\�|�������7�[��~�X��r%�q!eN�ҁF�Y(#h��'Mh��/>4<q����ޜ���ǔ�;�Ai�W�����8[���+��e�,�ǌj��(���t�ݏ�zn��A�\�(�x!,^�<�6����I�Y ��^r1dc������(~!�(3�"��L٨�L.I|"��׳��J��oY�N���'�O��<�V�Ss�<��[Z<��|7?���p�?�VA��Y��U�M�m�8���;�V/-D��-ysT�[�#��Z��9�䩗�1�?/��<�4K��Puj7�X�W����'����if##��D�u����t�KC�Q\��h� ���+N�9�x��G�G��é<��f����uto��aڿܬ_Z3��<��ϝO�5>K/ɟNjw8�%����L�~������[oړ3fJ�%���k������Q��x�53k��{ꐍ�{�������2bFC������K�� |��@�Ԧx�tz�>y�\�ƾ�<i� ����N�wt[�w/Q�{�X�-�-�uw��>�iv!8�w��}d�}9��w44�H��y:w��񛵍֐vC���aoK���dp%o�xq��:��l0����%Vf@����nN#\����׹��m�͓�ʜ2%�c�G|��|u8o���Lt�o��yT܆����|t���!��:Q�-\��l3�L�n<K{�]?`�o�_����a�=LǣҘ��i�t��{�G<U���x���4p����Q�$����7��iX�o�o�v �q��[��-<Ӹ�1K2� l?�0w�4��j���\�JM�8���/217�x����=�M*1a��<���
�ih�mo�j�g�9U�	t�3�-���y�o0�xRy� ���Kãr�a���_��N��(JGo̲TC��1D�0d�1�`��?A��e«8�f�x�[�.됭�ۺY�ao" �čf���6���?pO�G�f�V��Y,�4x�;:�������]<�58�Ec�L��m-���M��������?잺x
]��S ���E�2���WS�73�3��"�k����D!6�m򸔊���nqx���m�e9�t<�Ln$�h������͞��0�=�d�~�����#~�f&���ύ�:����h� Q�-e&����N^���HtC.n:6�Ã�6�k<�)~�i�4�5��۲��i��'�������R��&��Q���;4��?����.|�m���5O�	����`�?;:峇\�g��QC��Kޡ��������{�����kOSW�"�#/o���1����.ߙ�> Yӟ:#��F�mޖv3~�2���<��7�����v����o�]���[ou��5K�:���~½����������A���Q0�g�\4�of��h�Γ�K�ฃ�4M�X��`��T��6�������w��a���A8�o��yf}J.�HWZRO����q�JΧ�o�K�&��}��ʋQ��_�~:0w�����ɒC�b�[�x*<����z[}�v*�`�<�%����_�[��^���u {�[�]�iE��_�����h$r0e0ԷB@Q#�A�Ca�8��4s5m���r�ps����o�������t<��M�5����#����7=��v�=�o�֢�4�V��\��%@>���WaKF�����n:8?s?n���q���_M�ڞ6H��J����ˏ�ܴ���ছ}�g�W��V8;�$n��;�X��#�QA�?��y��#s#ms��w���VYs!�u��K�Ue�2R<NKJ���-�`k橐}��(�EcP�	�j��Z���O�?w͉Ϸ�w4tC�4�QF�<w��WI�*�9}x��a�[8\���a��y�m���sn�l�����7��F���H�%d>�G�����[�_&L�w���F��0:�M�A�����l&�`@�l�+Z�
=�����H��!;S��?�Z��A�U��!?���nw�N��ﹿ��l|!{���mO�*б�dvx�V���ձkح��V��`��`m�]���<a��a��d�Nr����mY�0�*p��c�9�����^��������Ki�dLaZ^W4^�;hK��_4�;�C�2��i:�a22\	��$nF�y���	����*ݍs�e��v��_�Lz6����Z1�~:\���ո۽��t�Cލû���h�Q�0��h[�xԯ`�[M��w(��q�]ş�v��k��e(����4i9����w�9�b>��;����v�p�;m_�7�MO{Lq�uo�����WS�1�ԔA1�!ǻ�=�4m�\�7\��p��'t'=K����i7ڶᕶUniw�s��##��C?b���<v�ٚ�CHv�r���<=�j��9����w(F�'w4-X|�isF�C̿�>ʬg|�{�7���w�턻���;�o美��f�
��;3_���h�ν���y�fF�C��mH�q���h'��0s�Xa<�0�>�_�c�0[�WÀ���v�c+��in���8=�>-+p�j+��u�鲢!W1��6p�����D��0��(a�6@�Uq���	��p�t�_\�Oƈ���dF����L�M�o:)�;Nx;mK^L������Mk�~��h�Ѯ���[�iK�:F�+��]�w�ѐ���I�?�QtH�?�JK���UK�s߀�t�7?M��M�}���ox����,{�Aӝ��� ���|�GX-[f��i��ɢ(3`*,�a�\w���u@�5�P��h(|h� �˸�|����ܷr�KL!3h�]�%/�a��e�iNǍ���)���
~;�Ig�G�AW�;�w?�I[�;�p_��Rɝoa�(��s�����w(�>�C�o\��m�o��<[2�|5B��1�fU�:��/@?�NH�e�ռ��w�H�0"���2�\���o⫙��I��������(?�Lì��_�F�'zSVoW턋Gj�2�$���%�;��y�a��g�*���š�s
=��?u�#�)�2���惡�<���*��}��It�1�+������~����������Q1��x���:�.�۱G�Q���Up�%c=�Ȩu�����4�m���c~��u��������0��z��
7���u���{�V�[	�<����8���ƺ��xޅ����q7���=�����l������q��o=�����_�m�/7���7N8���f�v9B����8��0d�F_0?���%L���5��Լj�VN���Ýi{�s�wn
~#�C��Ѱo12�>o��8����Έg;����3�wLˏY����lXv��G�����sƦe�Y)#06M+�Ï2����d{�J�/���U�	�Ė�s��j���Gӵry
~n��5�C��o#�#e�i���`w�{>*xw ����hR�:>��;��f�Jv��O��Z�S^P=��k���,>3f�����?J�O���Y��y g�u:��0�~�ૼŃ੎|��NeO�y�5NȚ�.K+�A��_㨎^q	��C�1KO�0�,��Po�³u�.���iC��7<�>e�:�}^'.���m: 4��˕�2x}�k��O�qj��g�rO���fm��7l&���zy�<�X)��V�FӴ�+����9�q󀽿�]��U�&}��,���7�j�7�7��m�������fc2h���U�m�#�B��I�:����^��լ��Vy�c�=d`���J�X���V��o����}�������������9��L_W��~#�^8�l�=n9��]v���Vj������=��o����w��f���{�������o�[���7s���;�x�tu��~�,na;|��]e�����������|���o}w��t�mZ�Ɯ�d�i�4�{�(�j&�ƽT��(׀xjyI��|�[}ڝ���-E�"_�f�W�S��� L��v]�V�t����?իh�45��G�tz{�5�Զ�O�6�t�c+]�������5[��@p5o� ��>�n�7�
Ұ�`ڒ��`U��|#����i<��Q}�B�x|��%�ӌ?�	��#)�<|�qt�¸����C-ejZ>�lűJ�*H�$e���R4�q�R��b�(K���1��,��ځ���[F>��u90-?�,����kԌUn�%�:%�	�t-��|)z������3q(<K���Wym|#�t$��2ʄ����/E�4�ָ����1p�[7.c\�WK�]�']?�N�2��#�
����W.sX�!��<!s��_��7�ܭݽ�4�s^�����i�6L�mFW������/c��҄�-�dc�I��{֟Mo���>h���t�c$/��s�m\�����wç�G��=����ܽ�;��˷��FK��(�Cu��E�6�u��y����̐��S���Tɩ2��uwNލ��MO�>��g}�7������?U|W<h�fh�poF|[��Ʒ*?#��?��ۉ�����    IEND�B`�PK   IqwT�/UK[  �     jsons/user_defined.json��Io�0��
�9��=ʭ-�P�BU�	�l�KB���	�J����̼�=O�1k	�$V�zm�cZ�P�	�� �/�֮U�r�9l���N�
��2�[���Bಜ�����s��)�y���)��$��_�I��U�u7E��2��Q�R�A7�I3D<����B�@��$��	Rn��1Ӳ��w��c�(¢�Rl;�����0�r�ă�0�ٻ�|�>�����f.�=�2�yPDIVx)�E�; �7�y
Շ��UN �t�����?]��o�����"�D�GĿ0�s��B��I%�z�����?/g�����e���~��η�PK   IqwTq�3B�  7f            ��    cirkitFile.jsonPK   IqwT�Ʈ�"^ /_ /           ��#  images/5007451c-e503-410b-b74d-3a3f8b63c8be.pngPK   IqwT�/UK[  �             ���u jsons/user_defined.jsonPK      �   "w   